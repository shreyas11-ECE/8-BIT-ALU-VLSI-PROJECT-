VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alu
  CLASS BLOCK ;
  FOREIGN alu ;
  ORIGIN 2.600 3.000 ;
  SIZE 156.400 BY 136.200 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 97.700 125.400 98.100 125.500 ;
        RECT 116.900 125.400 117.300 125.500 ;
        RECT 136.100 125.400 136.500 125.500 ;
        RECT 84.600 125.100 98.100 125.400 ;
        RECT 103.800 125.100 117.300 125.400 ;
        RECT 123.000 125.100 136.500 125.400 ;
        RECT 1.400 120.800 1.800 122.900 ;
        RECT 3.000 120.800 3.400 123.100 ;
        RECT 4.600 120.800 5.000 124.500 ;
        RECT 8.600 120.800 9.000 124.500 ;
        RECT 10.200 120.800 10.600 123.100 ;
        RECT 11.800 120.800 12.200 122.900 ;
        RECT 13.400 120.800 13.800 125.100 ;
        RECT 15.500 120.800 15.900 123.100 ;
        RECT 17.400 120.800 17.800 122.900 ;
        RECT 19.000 120.800 19.400 123.100 ;
        RECT 19.800 120.800 20.200 125.100 ;
        RECT 21.900 120.800 22.300 123.100 ;
        RECT 23.000 120.800 23.400 123.100 ;
        RECT 24.600 120.800 25.000 122.900 ;
        RECT 28.600 120.800 29.000 124.500 ;
        RECT 31.800 120.800 32.200 125.100 ;
        RECT 33.400 120.800 33.800 124.100 ;
        RECT 39.800 120.800 40.200 122.900 ;
        RECT 41.400 120.800 41.800 123.100 ;
        RECT 42.200 120.800 42.600 125.100 ;
        RECT 44.300 120.800 44.700 123.100 ;
        RECT 46.200 120.800 46.600 124.500 ;
        RECT 50.200 120.800 50.600 123.100 ;
        RECT 51.800 120.800 52.200 122.900 ;
        RECT 54.200 120.800 54.600 122.900 ;
        RECT 55.800 120.800 56.200 123.100 ;
        RECT 61.400 120.800 61.800 124.100 ;
        RECT 63.000 120.800 63.400 125.100 ;
        RECT 65.100 120.800 65.500 123.100 ;
        RECT 66.200 120.800 66.600 123.100 ;
        RECT 67.800 120.800 68.200 123.100 ;
        RECT 69.400 120.800 69.800 122.900 ;
        RECT 71.800 120.800 72.200 123.100 ;
        RECT 73.400 120.800 73.800 122.900 ;
        RECT 75.000 120.800 75.400 123.100 ;
        RECT 75.800 120.800 76.200 125.100 ;
        RECT 77.400 120.800 77.800 125.100 ;
        RECT 79.000 120.800 79.400 125.100 ;
        RECT 84.600 124.800 85.000 125.100 ;
        RECT 86.200 125.000 86.700 125.100 ;
        RECT 103.800 124.800 104.200 125.100 ;
        RECT 105.500 125.000 105.900 125.100 ;
        RECT 123.000 124.800 123.400 125.100 ;
        RECT 124.700 125.000 125.100 125.100 ;
        RECT 80.600 120.800 81.000 122.900 ;
        RECT 82.200 120.800 82.600 123.100 ;
        RECT 83.000 120.800 83.400 123.100 ;
        RECT 84.600 120.800 85.000 123.100 ;
        RECT 86.200 120.800 86.600 123.100 ;
        RECT 89.400 120.800 89.800 123.100 ;
        RECT 91.000 120.800 91.400 123.100 ;
        RECT 95.000 120.800 95.400 123.100 ;
        RECT 96.600 120.800 97.000 123.100 ;
        RECT 98.200 120.800 98.600 123.100 ;
        RECT 99.800 120.800 100.200 123.100 ;
        RECT 102.200 120.800 102.600 123.100 ;
        RECT 103.800 120.800 104.200 123.100 ;
        RECT 105.400 120.800 105.800 123.100 ;
        RECT 108.600 120.800 109.000 123.100 ;
        RECT 110.200 120.800 110.600 123.100 ;
        RECT 114.200 120.800 114.600 123.100 ;
        RECT 115.800 120.800 116.200 123.100 ;
        RECT 117.400 120.800 117.800 123.100 ;
        RECT 119.000 120.800 119.400 123.100 ;
        RECT 120.600 120.800 121.000 123.100 ;
        RECT 121.400 120.800 121.800 123.100 ;
        RECT 123.000 120.800 123.400 123.100 ;
        RECT 124.600 120.800 125.000 123.100 ;
        RECT 127.800 120.800 128.200 123.100 ;
        RECT 129.400 120.800 129.800 123.100 ;
        RECT 133.400 120.800 133.800 123.100 ;
        RECT 135.000 120.800 135.400 123.100 ;
        RECT 136.600 120.800 137.000 123.100 ;
        RECT 138.200 120.800 138.600 123.100 ;
        RECT 139.800 120.800 140.200 124.500 ;
        RECT 142.200 120.800 142.600 124.500 ;
        RECT 144.600 120.800 145.000 124.500 ;
        RECT 146.200 120.800 146.600 125.100 ;
        RECT 147.800 120.800 148.200 123.100 ;
        RECT 149.400 120.800 149.800 123.100 ;
        RECT 0.200 120.200 151.000 120.800 ;
        RECT 1.400 118.100 1.800 120.200 ;
        RECT 3.000 117.900 3.400 120.200 ;
        RECT 4.600 118.100 5.000 120.200 ;
        RECT 6.200 117.900 6.600 120.200 ;
        RECT 8.600 115.900 9.000 120.200 ;
        RECT 10.200 118.100 10.600 120.200 ;
        RECT 11.800 117.900 12.200 120.200 ;
        RECT 12.600 117.900 13.000 120.200 ;
        RECT 14.200 117.900 14.600 120.200 ;
        RECT 15.000 117.900 15.400 120.200 ;
        RECT 16.600 118.100 17.000 120.200 ;
        RECT 18.500 117.900 18.900 120.200 ;
        RECT 20.600 115.900 21.000 120.200 ;
        RECT 22.200 115.900 22.600 120.200 ;
        RECT 23.800 116.500 24.200 120.200 ;
        RECT 26.200 115.900 26.600 120.200 ;
        RECT 28.300 117.900 28.700 120.200 ;
        RECT 30.200 116.500 30.600 120.200 ;
        RECT 33.400 118.100 33.800 120.200 ;
        RECT 35.000 117.900 35.400 120.200 ;
        RECT 35.800 117.900 36.200 120.200 ;
        RECT 37.400 118.100 37.800 120.200 ;
        RECT 39.300 117.900 39.700 120.200 ;
        RECT 41.400 115.900 41.800 120.200 ;
        RECT 42.200 117.900 42.600 120.200 ;
        RECT 43.800 118.100 44.200 120.200 ;
        RECT 47.000 116.500 47.400 120.200 ;
        RECT 51.000 117.900 51.400 120.200 ;
        RECT 51.800 117.900 52.200 120.200 ;
        RECT 53.400 117.900 53.800 120.200 ;
        RECT 55.800 115.900 56.200 120.200 ;
        RECT 57.900 115.900 58.300 120.200 ;
        RECT 61.400 116.500 61.800 120.200 ;
        RECT 63.800 115.900 64.200 120.200 ;
        RECT 66.200 116.500 66.600 120.200 ;
        RECT 67.800 117.900 68.200 120.200 ;
        RECT 69.400 118.100 69.800 120.200 ;
        RECT 71.000 115.900 71.400 120.200 ;
        RECT 73.100 117.900 73.500 120.200 ;
        RECT 75.000 118.100 75.400 120.200 ;
        RECT 76.600 117.900 77.000 120.200 ;
        RECT 77.400 117.900 77.800 120.200 ;
        RECT 79.000 115.900 79.400 120.200 ;
        RECT 81.100 117.900 81.500 120.200 ;
        RECT 82.200 117.900 82.600 120.200 ;
        RECT 83.800 117.900 84.200 120.200 ;
        RECT 85.400 117.900 85.800 120.200 ;
        RECT 88.600 117.900 89.000 120.200 ;
        RECT 90.200 117.900 90.600 120.200 ;
        RECT 94.200 117.900 94.600 120.200 ;
        RECT 95.800 117.900 96.200 120.200 ;
        RECT 97.400 117.900 97.800 120.200 ;
        RECT 99.000 117.900 99.400 120.200 ;
        RECT 83.800 115.900 84.200 116.200 ;
        RECT 85.500 115.900 85.900 116.000 ;
        RECT 103.000 115.900 103.400 120.200 ;
        RECT 103.800 115.900 104.200 120.200 ;
        RECT 107.800 116.500 108.200 120.200 ;
        RECT 110.200 118.100 110.600 120.200 ;
        RECT 111.800 117.900 112.200 120.200 ;
        RECT 113.400 117.900 113.800 120.200 ;
        RECT 115.000 116.500 115.400 120.200 ;
        RECT 119.000 116.500 119.400 120.200 ;
        RECT 122.200 117.900 122.600 120.200 ;
        RECT 123.800 117.900 124.200 120.200 ;
        RECT 125.400 117.900 125.800 120.200 ;
        RECT 128.600 117.900 129.000 120.200 ;
        RECT 130.200 117.900 130.600 120.200 ;
        RECT 134.200 117.900 134.600 120.200 ;
        RECT 135.800 117.900 136.200 120.200 ;
        RECT 137.400 117.900 137.800 120.200 ;
        RECT 139.000 117.900 139.400 120.200 ;
        RECT 140.600 117.900 141.000 120.200 ;
        RECT 142.200 116.500 142.600 120.200 ;
        RECT 144.600 116.500 145.000 120.200 ;
        RECT 147.000 116.500 147.400 120.200 ;
        RECT 123.800 115.900 124.200 116.200 ;
        RECT 125.400 115.900 125.900 116.000 ;
        RECT 83.800 115.600 97.300 115.900 ;
        RECT 123.800 115.600 137.300 115.900 ;
        RECT 96.900 115.500 97.300 115.600 ;
        RECT 136.900 115.500 137.300 115.600 ;
        RECT 117.700 105.400 118.100 105.500 ;
        RECT 138.500 105.400 138.900 105.500 ;
        RECT 104.600 105.100 118.100 105.400 ;
        RECT 125.400 105.100 138.900 105.400 ;
        RECT 0.900 100.800 1.300 103.100 ;
        RECT 3.000 100.800 3.400 105.100 ;
        RECT 5.400 100.800 5.800 104.500 ;
        RECT 7.800 100.800 8.200 102.900 ;
        RECT 9.400 100.800 9.800 103.100 ;
        RECT 10.200 100.800 10.600 103.100 ;
        RECT 11.800 100.800 12.200 102.900 ;
        RECT 13.400 100.800 13.800 103.100 ;
        RECT 15.000 100.800 15.400 103.100 ;
        RECT 15.800 100.800 16.200 105.100 ;
        RECT 17.400 100.800 17.800 103.100 ;
        RECT 19.000 100.800 19.400 103.100 ;
        RECT 20.600 100.800 21.000 102.900 ;
        RECT 22.200 100.800 22.600 103.100 ;
        RECT 23.800 100.800 24.200 102.900 ;
        RECT 25.400 100.800 25.800 103.100 ;
        RECT 27.800 100.800 28.200 104.500 ;
        RECT 29.400 100.800 29.800 103.100 ;
        RECT 31.000 100.800 31.400 102.900 ;
        RECT 32.600 100.800 33.000 103.100 ;
        RECT 34.200 100.800 34.600 102.900 ;
        RECT 37.400 100.800 37.800 104.500 ;
        RECT 40.600 100.800 41.000 104.500 ;
        RECT 42.200 100.800 42.600 103.100 ;
        RECT 43.800 100.800 44.200 102.900 ;
        RECT 45.400 100.800 45.800 103.100 ;
        RECT 47.000 100.800 47.400 102.900 ;
        RECT 50.200 100.800 50.600 103.100 ;
        RECT 51.800 100.800 52.200 102.900 ;
        RECT 53.700 100.800 54.100 103.100 ;
        RECT 55.800 100.800 56.200 105.100 ;
        RECT 56.900 100.800 57.300 103.100 ;
        RECT 59.000 100.800 59.400 105.100 ;
        RECT 60.600 100.800 61.000 104.500 ;
        RECT 63.000 100.800 63.400 105.100 ;
        RECT 65.100 100.800 65.500 103.100 ;
        RECT 66.500 100.800 66.900 103.100 ;
        RECT 68.600 100.800 69.000 105.100 ;
        RECT 70.200 100.800 70.600 102.900 ;
        RECT 71.800 100.800 72.200 103.100 ;
        RECT 74.200 100.800 74.600 104.500 ;
        RECT 75.800 100.800 76.200 103.100 ;
        RECT 77.400 100.800 77.800 103.100 ;
        RECT 79.000 100.800 79.400 103.100 ;
        RECT 81.400 100.800 81.800 104.500 ;
        RECT 83.000 100.800 83.400 103.100 ;
        RECT 84.600 100.800 85.000 102.900 ;
        RECT 86.200 100.800 86.600 103.100 ;
        RECT 88.600 100.800 89.000 104.500 ;
        RECT 91.800 100.800 92.200 104.500 ;
        RECT 95.800 100.800 96.200 105.100 ;
        RECT 98.200 100.800 98.600 105.100 ;
        RECT 99.000 100.800 99.400 105.100 ;
        RECT 104.600 104.800 105.000 105.100 ;
        RECT 106.200 105.000 106.700 105.100 ;
        RECT 103.000 100.800 103.400 103.100 ;
        RECT 104.600 100.800 105.000 103.100 ;
        RECT 106.200 100.800 106.600 103.100 ;
        RECT 109.400 100.800 109.800 103.100 ;
        RECT 111.000 100.800 111.400 103.100 ;
        RECT 115.000 100.800 115.400 103.100 ;
        RECT 116.600 100.800 117.000 103.100 ;
        RECT 118.200 100.800 118.600 103.100 ;
        RECT 119.800 100.800 120.200 103.100 ;
        RECT 120.900 100.800 121.300 103.100 ;
        RECT 123.000 100.800 123.400 105.100 ;
        RECT 125.400 104.800 125.800 105.100 ;
        RECT 127.100 105.000 127.500 105.100 ;
        RECT 123.800 100.800 124.200 103.100 ;
        RECT 125.400 100.800 125.800 103.100 ;
        RECT 127.000 100.800 127.400 103.100 ;
        RECT 130.200 100.800 130.600 103.100 ;
        RECT 131.800 100.800 132.200 103.100 ;
        RECT 135.800 100.800 136.200 103.100 ;
        RECT 137.400 100.800 137.800 103.100 ;
        RECT 139.000 100.800 139.400 103.100 ;
        RECT 140.600 100.800 141.000 103.100 ;
        RECT 141.400 100.800 141.800 103.100 ;
        RECT 143.000 100.800 143.400 103.100 ;
        RECT 144.600 100.800 145.000 102.900 ;
        RECT 146.200 100.800 146.600 105.100 ;
        RECT 0.200 100.200 151.000 100.800 ;
        RECT 1.400 98.100 1.800 100.200 ;
        RECT 3.000 97.900 3.400 100.200 ;
        RECT 3.800 95.900 4.200 100.200 ;
        RECT 6.200 98.100 6.600 100.200 ;
        RECT 7.800 97.900 8.200 100.200 ;
        RECT 8.600 97.900 9.000 100.200 ;
        RECT 10.200 97.900 10.600 100.200 ;
        RECT 11.800 96.500 12.200 100.200 ;
        RECT 15.800 98.100 16.200 100.200 ;
        RECT 17.400 97.900 17.800 100.200 ;
        RECT 19.000 96.500 19.400 100.200 ;
        RECT 21.400 95.900 21.800 100.200 ;
        RECT 23.500 97.900 23.900 100.200 ;
        RECT 26.200 96.500 26.600 100.200 ;
        RECT 28.600 98.100 29.000 100.200 ;
        RECT 30.200 97.900 30.600 100.200 ;
        RECT 31.800 98.100 32.200 100.200 ;
        RECT 33.400 97.900 33.800 100.200 ;
        RECT 35.800 96.500 36.200 100.200 ;
        RECT 37.400 97.900 37.800 100.200 ;
        RECT 39.000 98.100 39.400 100.200 ;
        RECT 41.400 95.900 41.800 100.200 ;
        RECT 42.200 97.900 42.600 100.200 ;
        RECT 43.800 98.100 44.200 100.200 ;
        RECT 45.400 97.900 45.800 100.200 ;
        RECT 47.000 98.100 47.400 100.200 ;
        RECT 50.200 97.900 50.600 100.200 ;
        RECT 51.800 98.100 52.200 100.200 ;
        RECT 53.400 97.900 53.800 100.200 ;
        RECT 55.000 98.100 55.400 100.200 ;
        RECT 58.200 95.900 58.600 100.200 ;
        RECT 59.800 98.100 60.200 100.200 ;
        RECT 61.400 97.900 61.800 100.200 ;
        RECT 63.800 96.500 64.200 100.200 ;
        RECT 67.000 96.500 67.400 100.200 ;
        RECT 68.600 97.900 69.000 100.200 ;
        RECT 70.200 98.100 70.600 100.200 ;
        RECT 73.400 96.500 73.800 100.200 ;
        RECT 76.600 95.900 77.000 100.200 ;
        RECT 77.400 95.900 77.800 100.200 ;
        RECT 80.600 95.900 81.000 100.200 ;
        RECT 81.700 97.900 82.100 100.200 ;
        RECT 83.800 95.900 84.200 100.200 ;
        RECT 84.600 95.900 85.000 100.200 ;
        RECT 86.700 97.900 87.100 100.200 ;
        RECT 88.600 95.900 89.000 100.200 ;
        RECT 89.700 97.900 90.100 100.200 ;
        RECT 91.800 95.900 92.200 100.200 ;
        RECT 94.200 95.900 94.600 100.200 ;
        RECT 95.800 98.100 96.200 100.200 ;
        RECT 97.400 97.900 97.800 100.200 ;
        RECT 98.200 95.900 98.600 100.200 ;
        RECT 100.300 97.900 100.700 100.200 ;
        RECT 103.000 95.900 103.400 100.200 ;
        RECT 105.100 97.900 105.500 100.200 ;
        RECT 107.000 97.900 107.400 100.200 ;
        RECT 109.400 95.900 109.800 100.200 ;
        RECT 111.800 95.900 112.200 100.200 ;
        RECT 112.600 97.900 113.000 100.200 ;
        RECT 114.200 97.900 114.600 100.200 ;
        RECT 115.000 95.900 115.400 100.200 ;
        RECT 117.100 97.900 117.500 100.200 ;
        RECT 119.000 96.500 119.400 100.200 ;
        RECT 121.400 95.900 121.800 100.200 ;
        RECT 123.800 97.900 124.200 100.200 ;
        RECT 125.400 97.900 125.800 100.200 ;
        RECT 127.000 97.900 127.400 100.200 ;
        RECT 130.200 97.900 130.600 100.200 ;
        RECT 131.800 97.900 132.200 100.200 ;
        RECT 135.800 97.900 136.200 100.200 ;
        RECT 137.400 97.900 137.800 100.200 ;
        RECT 139.000 97.900 139.400 100.200 ;
        RECT 140.600 97.900 141.000 100.200 ;
        RECT 142.200 96.500 142.600 100.200 ;
        RECT 125.400 95.900 125.800 96.200 ;
        RECT 127.100 95.900 127.500 96.000 ;
        RECT 143.800 95.900 144.200 100.200 ;
        RECT 147.000 96.500 147.400 100.200 ;
        RECT 148.600 97.900 149.000 100.200 ;
        RECT 125.400 95.600 138.900 95.900 ;
        RECT 138.500 95.500 138.900 95.600 ;
        RECT 1.400 80.800 1.800 84.500 ;
        RECT 4.100 80.800 4.500 83.100 ;
        RECT 6.200 80.800 6.600 85.100 ;
        RECT 7.800 80.800 8.200 82.900 ;
        RECT 9.400 80.800 9.800 83.100 ;
        RECT 11.800 80.800 12.200 84.500 ;
        RECT 14.200 80.800 14.600 82.900 ;
        RECT 15.800 80.800 16.200 83.100 ;
        RECT 16.600 80.800 17.000 83.100 ;
        RECT 18.200 80.800 18.600 82.900 ;
        RECT 20.600 81.100 21.100 84.400 ;
        RECT 20.700 80.800 21.100 81.100 ;
        RECT 23.700 80.800 24.200 84.400 ;
        RECT 25.400 80.800 25.800 83.100 ;
        RECT 27.000 80.800 27.400 83.100 ;
        RECT 28.100 80.800 28.500 83.100 ;
        RECT 30.200 80.800 30.600 85.100 ;
        RECT 31.300 80.800 31.700 83.100 ;
        RECT 33.400 80.800 33.800 85.100 ;
        RECT 35.000 80.800 35.400 82.900 ;
        RECT 36.600 80.800 37.000 83.100 ;
        RECT 39.000 80.800 39.400 84.500 ;
        RECT 40.600 80.800 41.000 83.100 ;
        RECT 42.200 80.800 42.600 83.100 ;
        RECT 43.000 80.800 43.400 83.100 ;
        RECT 44.600 80.800 45.000 83.100 ;
        RECT 45.700 80.800 46.100 83.100 ;
        RECT 47.800 80.800 48.200 85.100 ;
        RECT 50.200 80.800 50.600 83.100 ;
        RECT 51.800 80.800 52.200 83.100 ;
        RECT 52.600 80.800 53.000 85.100 ;
        RECT 54.700 80.800 55.100 83.100 ;
        RECT 56.600 80.800 57.000 84.500 ;
        RECT 59.000 80.800 59.400 83.100 ;
        RECT 60.600 80.800 61.000 83.100 ;
        RECT 61.400 80.800 61.800 83.100 ;
        RECT 63.000 80.800 63.400 83.100 ;
        RECT 64.100 80.800 64.500 83.100 ;
        RECT 66.200 80.800 66.600 85.100 ;
        RECT 67.300 80.800 67.700 83.100 ;
        RECT 69.400 80.800 69.800 85.100 ;
        RECT 70.200 80.800 70.600 85.100 ;
        RECT 72.300 80.800 72.700 83.100 ;
        RECT 73.400 80.800 73.800 83.100 ;
        RECT 75.000 80.800 75.400 83.100 ;
        RECT 76.600 80.800 77.100 84.400 ;
        RECT 79.700 81.100 80.200 84.400 ;
        RECT 79.700 80.800 80.100 81.100 ;
        RECT 81.400 80.800 81.800 83.100 ;
        RECT 83.000 80.800 83.400 84.900 ;
        RECT 85.400 80.800 85.800 85.100 ;
        RECT 86.200 80.800 86.600 85.100 ;
        RECT 87.800 80.800 88.200 85.100 ;
        RECT 88.600 80.800 89.000 85.100 ;
        RECT 90.700 80.800 91.100 83.100 ;
        RECT 93.400 80.800 93.800 84.500 ;
        RECT 95.000 80.800 95.400 85.100 ;
        RECT 97.400 80.800 97.800 83.100 ;
        RECT 101.400 80.800 101.900 84.400 ;
        RECT 104.500 81.100 105.000 84.400 ;
        RECT 104.500 80.800 104.900 81.100 ;
        RECT 106.200 80.800 106.600 83.100 ;
        RECT 107.800 80.800 108.200 83.100 ;
        RECT 108.600 80.800 109.000 85.100 ;
        RECT 110.200 80.800 110.600 85.100 ;
        RECT 111.800 80.800 112.200 84.500 ;
        RECT 114.500 80.800 114.900 83.100 ;
        RECT 116.600 80.800 117.000 85.100 ;
        RECT 119.000 80.800 119.400 85.100 ;
        RECT 121.100 80.800 121.500 85.100 ;
        RECT 123.800 80.800 124.200 84.500 ;
        RECT 126.200 80.800 126.600 85.100 ;
        RECT 128.300 80.800 128.700 83.100 ;
        RECT 129.400 80.800 129.800 85.100 ;
        RECT 131.500 80.800 131.900 83.100 ;
        RECT 133.400 81.100 133.900 84.400 ;
        RECT 133.500 80.800 133.900 81.100 ;
        RECT 136.500 80.800 137.000 84.400 ;
        RECT 139.000 80.800 139.400 84.500 ;
        RECT 141.700 80.800 142.100 83.100 ;
        RECT 143.800 80.800 144.200 85.100 ;
        RECT 145.400 80.800 145.800 83.100 ;
        RECT 147.000 80.800 147.400 84.500 ;
        RECT 148.600 80.800 149.000 83.100 ;
        RECT 150.200 80.800 150.600 83.100 ;
        RECT 0.200 80.200 151.000 80.800 ;
        RECT 1.400 78.100 1.800 80.200 ;
        RECT 3.000 77.900 3.400 80.200 ;
        RECT 4.100 77.900 4.500 80.200 ;
        RECT 6.200 75.900 6.600 80.200 ;
        RECT 7.800 78.100 8.200 80.200 ;
        RECT 9.400 77.900 9.800 80.200 ;
        RECT 11.800 76.500 12.200 80.200 ;
        RECT 13.400 77.900 13.800 80.200 ;
        RECT 15.000 78.100 15.400 80.200 ;
        RECT 16.600 77.900 17.000 80.200 ;
        RECT 18.200 77.900 18.600 80.200 ;
        RECT 19.000 75.900 19.400 80.200 ;
        RECT 21.100 77.900 21.500 80.200 ;
        RECT 22.200 75.900 22.600 80.200 ;
        RECT 24.300 77.900 24.700 80.200 ;
        RECT 25.400 77.900 25.800 80.200 ;
        RECT 27.000 77.900 27.400 80.200 ;
        RECT 27.800 77.900 28.200 80.200 ;
        RECT 29.700 77.900 30.100 80.200 ;
        RECT 31.800 75.900 32.200 80.200 ;
        RECT 32.600 75.900 33.000 80.200 ;
        RECT 34.700 77.900 35.100 80.200 ;
        RECT 35.800 77.900 36.200 80.200 ;
        RECT 37.400 77.900 37.800 80.200 ;
        RECT 39.800 76.500 40.200 80.200 ;
        RECT 42.200 78.100 42.600 80.200 ;
        RECT 43.800 77.900 44.200 80.200 ;
        RECT 46.200 76.500 46.600 80.200 ;
        RECT 49.400 77.900 49.800 80.200 ;
        RECT 51.000 78.100 51.400 80.200 ;
        RECT 53.400 77.900 53.800 80.200 ;
        RECT 54.200 77.900 54.600 80.200 ;
        RECT 55.800 78.100 56.200 80.200 ;
        RECT 57.400 77.900 57.800 80.200 ;
        RECT 59.000 78.100 59.400 80.200 ;
        RECT 62.200 75.900 62.600 80.200 ;
        RECT 63.300 77.900 63.700 80.200 ;
        RECT 65.400 75.900 65.800 80.200 ;
        RECT 66.200 75.900 66.600 80.200 ;
        RECT 68.300 77.900 68.700 80.200 ;
        RECT 69.400 75.900 69.800 80.200 ;
        RECT 71.800 75.900 72.200 80.200 ;
        RECT 73.900 77.900 74.300 80.200 ;
        RECT 75.000 75.900 75.400 80.200 ;
        RECT 76.600 77.900 77.000 80.200 ;
        RECT 78.200 77.900 78.600 80.200 ;
        RECT 79.000 75.900 79.400 80.200 ;
        RECT 80.600 75.900 81.000 80.200 ;
        RECT 81.400 77.900 81.800 80.200 ;
        RECT 83.000 77.900 83.400 80.200 ;
        RECT 83.800 75.900 84.200 80.200 ;
        RECT 85.900 77.900 86.300 80.200 ;
        RECT 88.600 75.900 89.000 80.200 ;
        RECT 89.400 75.900 89.800 80.200 ;
        RECT 91.500 77.900 91.900 80.200 ;
        RECT 92.600 77.900 93.000 80.200 ;
        RECT 94.200 77.900 94.600 80.200 ;
        RECT 95.000 77.900 95.400 80.200 ;
        RECT 96.600 76.100 97.000 80.200 ;
        RECT 100.600 76.500 101.000 80.200 ;
        RECT 104.600 77.900 105.000 80.200 ;
        RECT 107.000 76.500 107.400 80.200 ;
        RECT 109.400 76.500 109.800 80.200 ;
        RECT 112.600 76.100 113.000 80.200 ;
        RECT 114.200 77.900 114.600 80.200 ;
        RECT 116.600 75.900 117.000 80.200 ;
        RECT 117.700 77.900 118.100 80.200 ;
        RECT 119.800 75.900 120.200 80.200 ;
        RECT 120.600 77.900 121.000 80.200 ;
        RECT 122.200 77.900 122.600 80.200 ;
        RECT 124.600 76.500 125.000 80.200 ;
        RECT 126.200 77.900 126.600 80.200 ;
        RECT 127.800 76.100 128.200 80.200 ;
        RECT 131.000 75.900 131.400 80.200 ;
        RECT 131.800 75.900 132.200 80.200 ;
        RECT 133.400 75.900 133.800 80.200 ;
        RECT 135.500 77.900 135.900 80.200 ;
        RECT 136.600 75.900 137.000 80.200 ;
        RECT 138.700 77.900 139.100 80.200 ;
        RECT 140.100 77.900 140.500 80.200 ;
        RECT 142.200 75.900 142.600 80.200 ;
        RECT 144.300 75.900 144.700 80.200 ;
        RECT 147.000 75.900 147.400 80.200 ;
        RECT 147.800 77.900 148.200 80.200 ;
        RECT 149.400 77.900 149.800 80.200 ;
        RECT 1.400 60.800 1.800 64.500 ;
        RECT 3.800 60.800 4.200 65.100 ;
        RECT 7.800 60.800 8.200 64.500 ;
        RECT 9.400 60.800 9.800 63.100 ;
        RECT 11.000 60.800 11.400 62.900 ;
        RECT 13.400 60.800 13.800 62.900 ;
        RECT 15.000 60.800 15.400 63.100 ;
        RECT 15.800 60.800 16.200 63.100 ;
        RECT 17.400 60.800 17.800 62.900 ;
        RECT 19.800 60.800 20.200 64.900 ;
        RECT 21.400 60.800 21.800 63.100 ;
        RECT 23.800 60.800 24.200 65.100 ;
        RECT 24.600 60.800 25.000 65.100 ;
        RECT 27.800 60.800 28.200 65.100 ;
        RECT 28.600 60.800 29.000 63.100 ;
        RECT 30.200 60.800 30.600 63.100 ;
        RECT 32.600 60.800 33.000 64.500 ;
        RECT 34.200 60.800 34.600 63.100 ;
        RECT 35.800 60.800 36.200 63.100 ;
        RECT 36.600 60.800 37.000 63.100 ;
        RECT 38.200 60.800 38.600 63.100 ;
        RECT 39.300 60.800 39.700 63.100 ;
        RECT 41.400 60.800 41.800 65.100 ;
        RECT 42.200 60.800 42.600 65.100 ;
        RECT 44.300 60.800 44.700 63.100 ;
        RECT 45.700 60.800 46.100 63.100 ;
        RECT 47.800 60.800 48.200 65.100 ;
        RECT 50.200 60.800 50.600 65.100 ;
        RECT 52.300 60.800 52.700 63.100 ;
        RECT 53.400 60.800 53.800 63.100 ;
        RECT 55.000 60.800 55.400 63.100 ;
        RECT 55.800 60.800 56.200 65.100 ;
        RECT 59.000 60.800 59.400 65.100 ;
        RECT 62.200 60.800 62.600 64.500 ;
        RECT 65.400 60.800 65.800 64.500 ;
        RECT 67.800 60.800 68.200 64.500 ;
        RECT 70.200 60.800 70.600 63.100 ;
        RECT 71.800 60.800 72.200 63.100 ;
        RECT 72.600 60.800 73.000 63.100 ;
        RECT 74.200 60.800 74.600 63.100 ;
        RECT 75.000 60.800 75.400 65.100 ;
        RECT 77.100 60.800 77.500 63.100 ;
        RECT 79.000 60.800 79.400 64.900 ;
        RECT 81.600 60.800 82.000 65.100 ;
        RECT 83.000 60.800 83.400 63.100 ;
        RECT 84.600 60.800 85.000 63.100 ;
        RECT 85.400 60.800 85.800 63.100 ;
        RECT 87.000 60.800 87.400 63.100 ;
        RECT 87.800 60.800 88.200 65.100 ;
        RECT 90.200 60.800 90.600 63.100 ;
        RECT 91.800 60.800 92.200 65.100 ;
        RECT 93.900 60.800 94.300 63.100 ;
        RECT 95.000 60.800 95.400 65.100 ;
        RECT 99.000 60.800 99.400 65.100 ;
        RECT 101.400 60.800 101.800 65.100 ;
        RECT 103.500 60.800 103.900 63.100 ;
        RECT 104.600 60.800 105.000 63.100 ;
        RECT 106.200 60.800 106.600 63.100 ;
        RECT 107.300 60.800 107.700 63.100 ;
        RECT 109.400 60.800 109.800 65.100 ;
        RECT 110.500 60.800 110.900 63.100 ;
        RECT 112.600 60.800 113.000 65.100 ;
        RECT 115.000 60.800 115.400 65.100 ;
        RECT 115.800 60.800 116.200 65.100 ;
        RECT 117.900 60.800 118.300 63.100 ;
        RECT 119.000 60.800 119.400 65.100 ;
        RECT 121.400 60.800 121.800 63.100 ;
        RECT 123.000 60.800 123.400 63.100 ;
        RECT 124.100 60.800 124.500 63.100 ;
        RECT 126.200 60.800 126.600 65.100 ;
        RECT 127.000 60.800 127.400 63.100 ;
        RECT 128.600 60.800 129.000 63.100 ;
        RECT 130.200 60.800 130.600 63.100 ;
        RECT 131.000 60.800 131.400 63.100 ;
        RECT 133.400 60.800 133.800 64.500 ;
        RECT 139.000 60.800 139.400 64.500 ;
        RECT 140.600 60.800 141.000 63.100 ;
        RECT 142.200 60.800 142.600 62.900 ;
        RECT 144.900 60.800 145.300 65.100 ;
        RECT 148.600 60.800 149.000 64.500 ;
        RECT 0.200 60.200 151.000 60.800 ;
        RECT 0.600 57.900 1.000 60.200 ;
        RECT 2.200 57.900 2.600 60.200 ;
        RECT 3.800 58.100 4.200 60.200 ;
        RECT 6.500 55.900 6.900 60.200 ;
        RECT 8.900 57.900 9.300 60.200 ;
        RECT 11.000 55.900 11.400 60.200 ;
        RECT 12.100 57.900 12.500 60.200 ;
        RECT 14.200 55.900 14.600 60.200 ;
        RECT 15.800 56.500 16.200 60.200 ;
        RECT 18.200 57.900 18.600 60.200 ;
        RECT 19.800 58.100 20.200 60.200 ;
        RECT 22.200 58.100 22.600 60.200 ;
        RECT 23.800 57.900 24.200 60.200 ;
        RECT 25.400 58.100 25.800 60.200 ;
        RECT 27.000 57.900 27.400 60.200 ;
        RECT 29.400 56.500 29.800 60.200 ;
        RECT 31.000 57.900 31.400 60.200 ;
        RECT 32.600 58.100 33.000 60.200 ;
        RECT 34.200 57.900 34.600 60.200 ;
        RECT 35.800 58.100 36.200 60.200 ;
        RECT 37.400 55.900 37.800 60.200 ;
        RECT 40.600 55.900 41.000 60.200 ;
        RECT 43.800 56.500 44.200 60.200 ;
        RECT 47.000 56.500 47.400 60.200 ;
        RECT 51.000 55.900 51.400 60.200 ;
        RECT 53.400 56.500 53.800 60.200 ;
        RECT 55.000 55.900 55.400 60.200 ;
        RECT 59.000 56.500 59.400 60.200 ;
        RECT 60.600 57.900 61.000 60.200 ;
        RECT 62.200 57.900 62.600 60.200 ;
        RECT 63.000 55.900 63.400 60.200 ;
        RECT 64.600 55.900 65.000 60.200 ;
        RECT 66.200 55.900 66.600 60.200 ;
        RECT 67.000 55.900 67.400 60.200 ;
        RECT 69.400 55.900 69.800 60.200 ;
        RECT 72.600 57.900 73.000 60.200 ;
        RECT 75.000 55.900 75.400 60.200 ;
        RECT 76.600 55.900 77.000 60.200 ;
        RECT 77.700 57.900 78.100 60.200 ;
        RECT 79.800 55.900 80.200 60.200 ;
        RECT 80.600 57.900 81.000 60.200 ;
        RECT 82.200 57.900 82.600 60.200 ;
        RECT 84.600 55.900 85.000 60.200 ;
        RECT 85.400 55.900 85.800 60.200 ;
        RECT 87.500 57.900 87.900 60.200 ;
        RECT 88.600 57.900 89.000 60.200 ;
        RECT 90.200 55.900 90.600 60.200 ;
        RECT 92.300 57.900 92.700 60.200 ;
        RECT 93.400 55.900 93.800 60.200 ;
        RECT 95.500 57.900 95.900 60.200 ;
        RECT 96.600 55.900 97.000 60.200 ;
        RECT 100.600 55.900 101.000 60.200 ;
        RECT 102.700 57.900 103.100 60.200 ;
        RECT 103.800 57.900 104.200 60.200 ;
        RECT 105.400 55.900 105.800 60.200 ;
        RECT 109.400 56.500 109.800 60.200 ;
        RECT 111.000 55.900 111.400 60.200 ;
        RECT 113.100 57.900 113.500 60.200 ;
        RECT 114.200 57.900 114.600 60.200 ;
        RECT 115.800 55.900 116.200 60.200 ;
        RECT 117.900 57.900 118.300 60.200 ;
        RECT 119.000 57.900 119.400 60.200 ;
        RECT 120.600 57.900 121.000 60.200 ;
        RECT 123.000 55.900 123.400 60.200 ;
        RECT 124.600 56.500 125.000 60.200 ;
        RECT 127.000 55.900 127.400 60.200 ;
        RECT 129.100 57.900 129.500 60.200 ;
        RECT 131.800 56.500 132.200 60.200 ;
        RECT 133.400 57.900 133.800 60.200 ;
        RECT 135.000 58.100 135.400 60.200 ;
        RECT 136.600 55.900 137.000 60.200 ;
        RECT 138.200 55.900 138.600 60.200 ;
        RECT 139.000 55.900 139.400 60.200 ;
        RECT 141.100 57.900 141.500 60.200 ;
        RECT 142.200 55.900 142.600 60.200 ;
        RECT 146.200 55.900 146.600 60.200 ;
        RECT 147.800 57.900 148.200 60.200 ;
        RECT 148.600 55.900 149.000 60.200 ;
        RECT 1.400 40.800 1.800 44.900 ;
        RECT 3.000 40.800 3.400 43.100 ;
        RECT 3.800 40.800 4.200 43.100 ;
        RECT 5.400 40.800 5.800 43.100 ;
        RECT 7.000 40.800 7.400 42.900 ;
        RECT 8.600 40.800 9.000 43.100 ;
        RECT 9.400 40.800 9.800 43.100 ;
        RECT 11.000 40.800 11.400 43.100 ;
        RECT 11.800 40.800 12.200 43.100 ;
        RECT 13.400 40.800 13.800 45.100 ;
        RECT 15.500 40.800 15.900 43.100 ;
        RECT 18.200 40.800 18.600 45.100 ;
        RECT 19.800 40.800 20.300 44.400 ;
        RECT 22.900 41.100 23.400 44.400 ;
        RECT 22.900 40.800 23.300 41.100 ;
        RECT 26.200 40.800 26.600 44.500 ;
        RECT 28.100 40.800 28.500 43.100 ;
        RECT 30.200 40.800 30.600 45.100 ;
        RECT 31.300 40.800 31.700 43.100 ;
        RECT 33.400 40.800 33.800 45.100 ;
        RECT 34.200 40.800 34.600 45.100 ;
        RECT 36.300 40.800 36.700 43.100 ;
        RECT 37.700 40.800 38.100 43.100 ;
        RECT 39.800 40.800 40.200 45.100 ;
        RECT 42.200 40.800 42.600 45.100 ;
        RECT 44.600 40.800 45.000 44.500 ;
        RECT 46.200 40.800 46.600 43.100 ;
        RECT 47.800 40.800 48.200 43.100 ;
        RECT 51.800 40.800 52.200 44.500 ;
        RECT 53.400 40.800 53.800 43.100 ;
        RECT 55.000 40.800 55.400 43.100 ;
        RECT 55.800 40.800 56.200 43.100 ;
        RECT 57.400 40.800 57.800 43.100 ;
        RECT 58.500 40.800 58.900 43.100 ;
        RECT 60.600 40.800 61.000 45.100 ;
        RECT 61.400 40.800 61.800 43.100 ;
        RECT 63.000 40.800 63.400 43.100 ;
        RECT 63.800 40.800 64.200 45.100 ;
        RECT 65.400 40.800 65.800 44.500 ;
        RECT 67.800 40.800 68.200 44.500 ;
        RECT 69.400 40.800 69.800 45.100 ;
        RECT 70.200 40.800 70.600 43.100 ;
        RECT 71.800 40.800 72.200 43.100 ;
        RECT 72.600 40.800 73.000 43.100 ;
        RECT 74.200 40.800 74.600 43.100 ;
        RECT 75.300 40.800 75.700 43.100 ;
        RECT 77.400 40.800 77.800 45.100 ;
        RECT 79.800 40.800 80.200 45.100 ;
        RECT 80.600 40.800 81.000 45.100 ;
        RECT 82.700 40.800 83.100 43.100 ;
        RECT 83.800 40.800 84.200 45.100 ;
        RECT 85.900 40.800 86.300 43.100 ;
        RECT 87.300 40.800 87.700 43.100 ;
        RECT 89.400 40.800 89.800 45.100 ;
        RECT 90.200 40.800 90.600 45.100 ;
        RECT 92.300 40.800 92.700 43.100 ;
        RECT 93.400 40.800 93.800 43.100 ;
        RECT 95.000 40.800 95.400 43.100 ;
        RECT 95.800 40.800 96.200 45.100 ;
        RECT 97.900 40.800 98.300 43.100 ;
        RECT 100.600 40.800 101.000 45.100 ;
        RECT 103.800 40.800 104.200 45.100 ;
        RECT 104.900 40.800 105.300 43.100 ;
        RECT 107.000 40.800 107.400 45.100 ;
        RECT 107.800 40.800 108.200 45.100 ;
        RECT 109.900 40.800 110.300 43.100 ;
        RECT 111.800 40.800 112.200 43.100 ;
        RECT 112.600 40.800 113.000 45.100 ;
        RECT 115.000 40.800 115.400 45.100 ;
        RECT 117.100 40.800 117.500 43.100 ;
        RECT 118.200 40.800 118.600 45.100 ;
        RECT 120.300 40.800 120.700 43.100 ;
        RECT 121.400 40.800 121.800 43.100 ;
        RECT 123.000 40.800 123.400 43.100 ;
        RECT 124.600 40.800 125.000 44.500 ;
        RECT 127.300 40.800 127.700 43.100 ;
        RECT 129.400 40.800 129.800 45.100 ;
        RECT 130.200 40.800 130.600 43.100 ;
        RECT 131.800 40.800 132.200 42.900 ;
        RECT 134.200 40.800 134.600 45.100 ;
        RECT 135.000 40.800 135.400 45.100 ;
        RECT 137.400 40.800 137.800 45.100 ;
        RECT 139.000 40.800 139.400 45.100 ;
        RECT 140.600 40.800 141.000 44.500 ;
        RECT 143.000 40.800 143.400 43.100 ;
        RECT 144.600 40.800 145.000 43.100 ;
        RECT 145.700 40.800 146.100 43.100 ;
        RECT 147.800 40.800 148.200 45.100 ;
        RECT 148.600 40.800 149.000 45.100 ;
        RECT 0.200 40.200 151.000 40.800 ;
        RECT 0.900 37.900 1.300 40.200 ;
        RECT 3.000 35.900 3.400 40.200 ;
        RECT 4.600 36.500 5.000 40.200 ;
        RECT 7.000 37.900 7.400 40.200 ;
        RECT 8.600 38.100 9.000 40.200 ;
        RECT 10.200 35.900 10.600 40.200 ;
        RECT 12.300 37.900 12.700 40.200 ;
        RECT 13.400 37.900 13.800 40.200 ;
        RECT 15.000 38.100 15.400 40.200 ;
        RECT 18.200 36.500 18.600 40.200 ;
        RECT 19.800 37.900 20.200 40.200 ;
        RECT 21.400 38.100 21.800 40.200 ;
        RECT 23.900 39.900 24.300 40.200 ;
        RECT 23.800 36.600 24.300 39.900 ;
        RECT 26.900 36.600 27.400 40.200 ;
        RECT 28.600 37.900 29.000 40.200 ;
        RECT 30.200 37.900 30.600 40.200 ;
        RECT 31.800 37.900 32.200 40.200 ;
        RECT 33.400 36.500 33.800 40.200 ;
        RECT 35.000 35.900 35.400 40.200 ;
        RECT 35.800 37.900 36.200 40.200 ;
        RECT 37.400 37.900 37.800 40.200 ;
        RECT 39.000 36.500 39.400 40.200 ;
        RECT 40.600 35.900 41.000 40.200 ;
        RECT 43.800 36.500 44.200 40.200 ;
        RECT 45.400 37.900 45.800 40.200 ;
        RECT 47.000 37.900 47.400 40.200 ;
        RECT 49.400 35.900 49.800 40.200 ;
        RECT 51.000 36.500 51.400 40.200 ;
        RECT 53.400 36.500 53.800 40.200 ;
        RECT 55.000 35.900 55.400 40.200 ;
        RECT 56.600 36.500 57.000 40.200 ;
        RECT 58.200 35.900 58.600 40.200 ;
        RECT 59.800 36.100 60.200 40.200 ;
        RECT 62.400 35.900 62.800 40.200 ;
        RECT 64.400 35.900 64.800 40.200 ;
        RECT 67.000 36.100 67.400 40.200 ;
        RECT 68.600 35.900 69.000 40.200 ;
        RECT 70.700 37.900 71.100 40.200 ;
        RECT 72.600 36.500 73.000 40.200 ;
        RECT 75.000 35.900 75.400 40.200 ;
        RECT 77.100 37.900 77.500 40.200 ;
        RECT 78.500 37.900 78.900 40.200 ;
        RECT 80.600 35.900 81.000 40.200 ;
        RECT 81.400 35.900 81.800 40.200 ;
        RECT 83.500 37.900 83.900 40.200 ;
        RECT 84.600 37.900 85.000 40.200 ;
        RECT 86.200 37.900 86.600 40.200 ;
        RECT 87.000 35.900 87.400 40.200 ;
        RECT 91.000 36.500 91.400 40.200 ;
        RECT 94.200 35.900 94.600 40.200 ;
        RECT 95.000 35.900 95.400 40.200 ;
        RECT 97.100 37.900 97.500 40.200 ;
        RECT 99.800 36.500 100.200 40.200 ;
        RECT 103.000 37.900 103.400 40.200 ;
        RECT 104.600 37.900 105.000 40.200 ;
        RECT 106.200 35.900 106.600 40.200 ;
        RECT 107.300 37.900 107.700 40.200 ;
        RECT 109.400 35.900 109.800 40.200 ;
        RECT 111.800 35.900 112.200 40.200 ;
        RECT 112.600 37.900 113.000 40.200 ;
        RECT 114.200 36.100 114.600 40.200 ;
        RECT 115.800 35.900 116.200 40.200 ;
        RECT 117.900 37.900 118.300 40.200 ;
        RECT 119.000 37.900 119.400 40.200 ;
        RECT 120.600 37.900 121.000 40.200 ;
        RECT 122.700 35.900 123.100 40.200 ;
        RECT 125.400 36.500 125.800 40.200 ;
        RECT 127.800 35.900 128.200 40.200 ;
        RECT 131.300 35.900 131.700 40.200 ;
        RECT 134.200 35.900 134.600 40.200 ;
        RECT 135.800 38.100 136.200 40.200 ;
        RECT 137.400 37.900 137.800 40.200 ;
        RECT 139.300 35.900 139.700 40.200 ;
        RECT 143.000 35.900 143.400 40.200 ;
        RECT 143.800 37.900 144.200 40.200 ;
        RECT 145.400 37.900 145.800 40.200 ;
        RECT 147.300 35.900 147.700 40.200 ;
        RECT 1.400 20.800 1.900 24.400 ;
        RECT 4.500 21.100 5.000 24.400 ;
        RECT 4.500 20.800 4.900 21.100 ;
        RECT 7.000 20.800 7.400 22.900 ;
        RECT 8.600 20.800 9.000 23.100 ;
        RECT 10.200 20.800 10.600 24.500 ;
        RECT 12.600 20.800 13.000 23.100 ;
        RECT 15.800 20.800 16.200 24.500 ;
        RECT 17.400 20.800 17.800 23.100 ;
        RECT 19.000 20.800 19.400 22.900 ;
        RECT 20.600 20.800 21.000 23.100 ;
        RECT 22.200 20.800 22.600 23.100 ;
        RECT 23.800 20.800 24.200 22.900 ;
        RECT 25.400 20.800 25.800 23.100 ;
        RECT 27.000 20.800 27.400 22.900 ;
        RECT 28.600 20.800 29.000 23.100 ;
        RECT 29.400 20.800 29.800 25.100 ;
        RECT 31.000 20.800 31.400 24.500 ;
        RECT 33.400 20.800 33.800 24.500 ;
        RECT 35.000 20.800 35.400 25.100 ;
        RECT 35.800 20.800 36.200 25.100 ;
        RECT 39.000 20.800 39.400 25.100 ;
        RECT 40.600 20.800 41.000 22.900 ;
        RECT 42.200 20.800 42.600 23.100 ;
        RECT 43.000 20.800 43.400 23.100 ;
        RECT 44.600 20.800 45.000 22.900 ;
        RECT 46.200 20.800 46.600 25.100 ;
        RECT 47.800 20.800 48.200 24.500 ;
        RECT 51.000 20.800 51.400 25.100 ;
        RECT 52.600 20.800 53.000 25.100 ;
        RECT 53.400 20.800 53.800 23.100 ;
        RECT 55.000 20.800 55.400 23.100 ;
        RECT 56.100 20.800 56.500 23.100 ;
        RECT 58.200 20.800 58.600 25.100 ;
        RECT 59.800 20.800 60.200 24.900 ;
        RECT 61.400 20.800 61.800 23.100 ;
        RECT 62.200 20.800 62.600 23.100 ;
        RECT 63.800 20.800 64.200 23.100 ;
        RECT 65.400 20.800 65.800 23.100 ;
        RECT 66.500 20.800 66.900 23.100 ;
        RECT 68.600 20.800 69.000 25.100 ;
        RECT 69.400 20.800 69.800 23.100 ;
        RECT 71.000 20.800 71.400 23.100 ;
        RECT 72.400 20.800 72.800 25.100 ;
        RECT 75.000 20.800 75.400 24.900 ;
        RECT 78.200 20.800 78.600 25.100 ;
        RECT 79.000 20.800 79.400 23.100 ;
        RECT 81.400 20.800 81.800 24.500 ;
        RECT 83.800 20.800 84.200 25.100 ;
        RECT 85.900 20.800 86.300 23.100 ;
        RECT 87.300 20.800 87.700 23.100 ;
        RECT 89.400 20.800 89.800 25.100 ;
        RECT 91.000 20.800 91.400 23.100 ;
        RECT 93.400 20.800 93.800 25.100 ;
        RECT 95.000 20.800 95.400 24.500 ;
        RECT 97.400 20.800 97.800 23.100 ;
        RECT 99.000 20.800 99.400 23.100 ;
        RECT 101.400 20.800 101.800 23.100 ;
        RECT 103.000 20.800 103.400 24.900 ;
        RECT 105.400 20.800 105.800 23.100 ;
        RECT 106.500 20.800 106.900 23.100 ;
        RECT 108.600 20.800 109.000 25.100 ;
        RECT 110.200 20.800 110.600 24.500 ;
        RECT 113.400 20.800 113.800 24.500 ;
        RECT 116.600 20.800 117.000 24.500 ;
        RECT 119.300 20.800 119.700 23.100 ;
        RECT 121.400 20.800 121.800 25.100 ;
        RECT 122.500 20.800 122.900 23.100 ;
        RECT 124.600 20.800 125.000 25.100 ;
        RECT 125.400 20.800 125.800 23.100 ;
        RECT 127.000 20.800 127.400 24.900 ;
        RECT 128.600 20.800 129.000 23.100 ;
        RECT 130.200 20.800 130.600 23.100 ;
        RECT 132.600 20.800 133.000 25.100 ;
        RECT 133.400 20.800 133.800 25.100 ;
        RECT 135.500 20.800 135.900 23.100 ;
        RECT 137.400 20.800 137.800 24.500 ;
        RECT 139.800 20.800 140.200 25.100 ;
        RECT 141.400 20.800 141.800 25.100 ;
        RECT 143.000 20.800 143.400 25.100 ;
        RECT 143.800 20.800 144.200 25.100 ;
        RECT 147.800 20.800 148.200 25.100 ;
        RECT 148.600 20.800 149.000 23.100 ;
        RECT 0.200 20.200 151.000 20.800 ;
        RECT 1.400 18.100 1.800 20.200 ;
        RECT 3.000 17.900 3.400 20.200 ;
        RECT 4.600 18.100 5.000 20.200 ;
        RECT 6.200 17.900 6.600 20.200 ;
        RECT 7.300 17.900 7.700 20.200 ;
        RECT 9.400 15.900 9.800 20.200 ;
        RECT 11.800 16.500 12.200 20.200 ;
        RECT 13.700 17.900 14.100 20.200 ;
        RECT 15.800 15.900 16.200 20.200 ;
        RECT 16.600 15.900 17.000 20.200 ;
        RECT 18.700 17.900 19.100 20.200 ;
        RECT 20.600 18.100 21.000 20.200 ;
        RECT 22.200 17.900 22.600 20.200 ;
        RECT 23.000 17.900 23.400 20.200 ;
        RECT 24.600 18.100 25.000 20.200 ;
        RECT 27.800 16.500 28.200 20.200 ;
        RECT 29.400 17.900 29.800 20.200 ;
        RECT 31.000 17.900 31.400 20.200 ;
        RECT 31.800 17.900 32.200 20.200 ;
        RECT 33.400 16.100 33.800 20.200 ;
        RECT 35.800 18.100 36.200 20.200 ;
        RECT 37.400 17.900 37.800 20.200 ;
        RECT 39.800 16.500 40.200 20.200 ;
        RECT 41.400 17.900 41.800 20.200 ;
        RECT 43.800 16.500 44.200 20.200 ;
        RECT 45.400 15.900 45.800 20.200 ;
        RECT 47.800 16.500 48.200 20.200 ;
        RECT 51.800 16.500 52.200 20.200 ;
        RECT 55.000 16.500 55.400 20.200 ;
        RECT 56.600 15.900 57.000 20.200 ;
        RECT 58.000 15.900 58.400 20.200 ;
        RECT 60.600 16.100 61.000 20.200 ;
        RECT 62.200 17.900 62.600 20.200 ;
        RECT 65.400 15.900 65.800 20.200 ;
        RECT 66.200 15.900 66.600 20.200 ;
        RECT 69.400 15.900 69.800 20.200 ;
        RECT 70.200 15.900 70.600 20.200 ;
        RECT 72.300 17.900 72.700 20.200 ;
        RECT 73.400 17.900 73.800 20.200 ;
        RECT 75.000 18.100 75.400 20.200 ;
        RECT 76.600 17.900 77.000 20.200 ;
        RECT 78.200 15.900 78.600 20.200 ;
        RECT 81.500 19.900 81.900 20.200 ;
        RECT 81.400 16.600 81.900 19.900 ;
        RECT 84.500 16.600 85.000 20.200 ;
        RECT 86.500 17.900 86.900 20.200 ;
        RECT 88.600 15.900 89.000 20.200 ;
        RECT 89.400 15.900 89.800 20.200 ;
        RECT 91.800 16.500 92.200 20.200 ;
        RECT 94.500 17.900 94.900 20.200 ;
        RECT 96.600 15.900 97.000 20.200 ;
        RECT 98.200 16.100 98.600 20.200 ;
        RECT 99.800 17.900 100.200 20.200 ;
        RECT 102.200 15.900 102.600 20.200 ;
        RECT 104.600 15.900 105.000 20.200 ;
        RECT 106.700 17.900 107.100 20.200 ;
        RECT 107.800 15.900 108.200 20.200 ;
        RECT 109.900 17.900 110.300 20.200 ;
        RECT 111.000 15.900 111.400 20.200 ;
        RECT 114.200 15.900 114.600 20.200 ;
        RECT 116.600 15.900 117.000 20.200 ;
        RECT 118.200 16.100 118.600 20.200 ;
        RECT 119.800 17.900 120.200 20.200 ;
        RECT 122.200 15.900 122.600 20.200 ;
        RECT 123.800 15.900 124.200 20.200 ;
        RECT 124.600 15.900 125.000 20.200 ;
        RECT 127.000 15.900 127.400 20.200 ;
        RECT 128.600 15.900 129.000 20.200 ;
        RECT 130.700 17.900 131.100 20.200 ;
        RECT 131.800 17.900 132.200 20.200 ;
        RECT 133.400 18.100 133.800 20.200 ;
        RECT 135.000 15.900 135.400 20.200 ;
        RECT 137.400 15.900 137.800 20.200 ;
        RECT 140.600 15.900 141.000 20.200 ;
        RECT 142.200 16.900 142.600 20.200 ;
        RECT 149.400 15.900 149.800 20.200 ;
        RECT 1.400 1.100 1.900 4.400 ;
        RECT 1.500 0.800 1.900 1.100 ;
        RECT 4.500 0.800 5.000 4.400 ;
        RECT 7.000 1.100 7.500 4.400 ;
        RECT 7.100 0.800 7.500 1.100 ;
        RECT 10.100 0.800 10.600 4.400 ;
        RECT 16.600 0.800 17.000 4.100 ;
        RECT 19.000 0.800 19.500 4.400 ;
        RECT 22.100 1.100 22.600 4.400 ;
        RECT 22.100 0.800 22.500 1.100 ;
        RECT 23.800 0.800 24.200 3.100 ;
        RECT 25.700 0.800 26.100 3.100 ;
        RECT 27.800 0.800 28.200 5.100 ;
        RECT 29.400 1.100 29.900 4.400 ;
        RECT 29.500 0.800 29.900 1.100 ;
        RECT 32.500 0.800 33.000 4.400 ;
        RECT 35.000 0.800 35.400 4.100 ;
        RECT 45.400 0.800 45.800 4.100 ;
        RECT 47.000 0.800 47.400 5.100 ;
        RECT 49.100 0.800 49.500 3.100 ;
        RECT 51.800 0.800 52.200 3.100 ;
        RECT 53.400 0.800 53.800 3.100 ;
        RECT 55.000 0.800 55.400 4.500 ;
        RECT 56.600 0.800 57.000 5.100 ;
        RECT 57.400 0.800 57.800 3.100 ;
        RECT 59.000 0.800 59.400 3.100 ;
        RECT 60.600 0.800 61.000 4.500 ;
        RECT 62.200 0.800 62.600 5.100 ;
        RECT 63.000 0.800 63.400 3.100 ;
        RECT 64.600 0.800 65.000 3.100 ;
        RECT 65.400 0.800 65.800 5.100 ;
        RECT 67.800 0.800 68.200 5.100 ;
        RECT 69.400 0.800 69.800 5.100 ;
        RECT 72.600 0.800 73.000 5.100 ;
        RECT 73.400 0.800 73.800 5.100 ;
        RECT 75.800 0.800 76.200 5.100 ;
        RECT 77.900 0.800 78.300 3.100 ;
        RECT 79.000 0.800 79.400 5.100 ;
        RECT 81.100 0.800 81.500 3.100 ;
        RECT 82.200 0.800 82.600 5.100 ;
        RECT 84.600 0.800 85.000 3.100 ;
        RECT 87.800 0.800 88.200 5.100 ;
        RECT 88.900 0.800 89.300 3.100 ;
        RECT 91.000 0.800 91.400 5.100 ;
        RECT 92.100 0.800 92.500 3.100 ;
        RECT 94.200 0.800 94.600 5.100 ;
        RECT 95.000 0.800 95.400 5.100 ;
        RECT 98.200 0.800 98.600 5.100 ;
        RECT 100.600 0.800 101.000 5.100 ;
        RECT 102.700 0.800 103.100 3.100 ;
        RECT 104.600 0.800 105.000 3.100 ;
        RECT 105.400 0.800 105.800 5.100 ;
        RECT 107.500 0.800 107.900 3.100 ;
        RECT 108.600 0.800 109.000 5.100 ;
        RECT 111.000 0.800 111.400 3.100 ;
        RECT 112.600 0.800 113.000 5.100 ;
        RECT 115.800 0.800 116.200 5.100 ;
        RECT 117.900 0.800 118.300 5.100 ;
        RECT 120.100 0.800 120.500 3.100 ;
        RECT 122.200 0.800 122.600 5.100 ;
        RECT 123.000 0.800 123.400 5.100 ;
        RECT 125.400 0.800 125.800 3.100 ;
        RECT 127.000 0.800 127.400 3.100 ;
        RECT 127.800 0.800 128.200 3.100 ;
        RECT 129.400 0.800 129.800 5.100 ;
        RECT 131.500 0.800 131.900 3.100 ;
        RECT 134.200 0.800 134.600 5.100 ;
        RECT 135.000 0.800 135.400 5.100 ;
        RECT 137.900 0.800 138.300 5.100 ;
        RECT 140.600 0.800 141.000 4.500 ;
        RECT 143.800 0.800 144.200 4.500 ;
        RECT 146.200 0.800 146.600 5.100 ;
        RECT 148.300 0.800 148.700 3.100 ;
        RECT 0.200 0.200 151.000 0.800 ;
      LAYER via1 ;
        RECT 86.200 122.700 86.600 123.100 ;
        RECT 103.800 121.800 104.200 122.200 ;
        RECT 123.000 121.800 123.400 122.200 ;
        RECT 48.200 120.300 48.600 120.700 ;
        RECT 48.900 120.300 49.300 120.700 ;
        RECT 83.800 118.800 84.200 119.200 ;
        RECT 83.800 115.800 84.200 116.200 ;
        RECT 125.400 118.800 125.800 119.200 ;
        RECT 125.400 115.600 125.800 116.000 ;
        RECT 106.200 102.700 106.600 103.100 ;
        RECT 125.400 101.800 125.800 102.200 ;
        RECT 48.200 100.300 48.600 100.700 ;
        RECT 48.900 100.300 49.300 100.700 ;
        RECT 125.400 98.800 125.800 99.200 ;
        RECT 125.400 95.800 125.800 96.200 ;
        RECT 48.200 80.300 48.600 80.700 ;
        RECT 48.900 80.300 49.300 80.700 ;
        RECT 48.200 60.300 48.600 60.700 ;
        RECT 48.900 60.300 49.300 60.700 ;
        RECT 48.200 40.300 48.600 40.700 ;
        RECT 48.900 40.300 49.300 40.700 ;
        RECT 48.200 20.300 48.600 20.700 ;
        RECT 48.900 20.300 49.300 20.700 ;
        RECT 48.200 0.300 48.600 0.700 ;
        RECT 48.900 0.300 49.300 0.700 ;
      LAYER metal2 ;
        RECT 86.200 125.000 86.600 125.400 ;
        RECT 86.200 123.100 86.500 125.000 ;
        RECT 103.800 124.800 104.200 125.200 ;
        RECT 123.000 124.800 123.400 125.200 ;
        RECT 86.200 122.700 86.600 123.100 ;
        RECT 103.800 122.200 104.100 124.800 ;
        RECT 123.000 122.200 123.300 124.800 ;
        RECT 103.800 121.800 104.200 122.200 ;
        RECT 123.000 121.800 123.400 122.200 ;
        RECT 48.000 120.300 49.600 120.700 ;
        RECT 83.800 118.800 84.200 119.200 ;
        RECT 125.400 118.800 125.800 119.200 ;
        RECT 83.800 116.200 84.100 118.800 ;
        RECT 83.800 115.800 84.200 116.200 ;
        RECT 125.400 116.000 125.700 118.800 ;
        RECT 125.400 115.600 125.800 116.000 ;
        RECT 106.200 105.000 106.600 105.400 ;
        RECT 106.200 103.100 106.500 105.000 ;
        RECT 125.400 104.800 125.800 105.200 ;
        RECT 106.200 102.700 106.600 103.100 ;
        RECT 125.400 102.200 125.700 104.800 ;
        RECT 125.400 101.800 125.800 102.200 ;
        RECT 48.000 100.300 49.600 100.700 ;
        RECT 125.400 98.800 125.800 99.200 ;
        RECT 125.400 96.200 125.700 98.800 ;
        RECT 125.400 95.800 125.800 96.200 ;
        RECT 48.000 80.300 49.600 80.700 ;
        RECT 48.000 60.300 49.600 60.700 ;
        RECT 48.000 40.300 49.600 40.700 ;
        RECT 48.000 20.300 49.600 20.700 ;
        RECT 48.000 0.300 49.600 0.700 ;
      LAYER via2 ;
        RECT 48.200 120.300 48.600 120.700 ;
        RECT 48.900 120.300 49.300 120.700 ;
        RECT 48.200 100.300 48.600 100.700 ;
        RECT 48.900 100.300 49.300 100.700 ;
        RECT 48.200 80.300 48.600 80.700 ;
        RECT 48.900 80.300 49.300 80.700 ;
        RECT 48.200 60.300 48.600 60.700 ;
        RECT 48.900 60.300 49.300 60.700 ;
        RECT 48.200 40.300 48.600 40.700 ;
        RECT 48.900 40.300 49.300 40.700 ;
        RECT 48.200 20.300 48.600 20.700 ;
        RECT 48.900 20.300 49.300 20.700 ;
        RECT 48.200 0.300 48.600 0.700 ;
        RECT 48.900 0.300 49.300 0.700 ;
      LAYER metal3 ;
        RECT 48.000 120.300 49.600 120.700 ;
        RECT 48.000 100.300 49.600 100.700 ;
        RECT 48.000 80.300 49.600 80.700 ;
        RECT 48.000 60.300 49.600 60.700 ;
        RECT 48.000 40.300 49.600 40.700 ;
        RECT 48.000 20.300 49.600 20.700 ;
        RECT 48.000 0.300 49.600 0.700 ;
      LAYER via3 ;
        RECT 48.200 120.300 48.600 120.700 ;
        RECT 49.000 120.300 49.400 120.700 ;
        RECT 48.200 100.300 48.600 100.700 ;
        RECT 49.000 100.300 49.400 100.700 ;
        RECT 48.200 80.300 48.600 80.700 ;
        RECT 49.000 80.300 49.400 80.700 ;
        RECT 48.200 60.300 48.600 60.700 ;
        RECT 49.000 60.300 49.400 60.700 ;
        RECT 48.200 40.300 48.600 40.700 ;
        RECT 49.000 40.300 49.400 40.700 ;
        RECT 48.200 20.300 48.600 20.700 ;
        RECT 49.000 20.300 49.400 20.700 ;
        RECT 48.200 0.300 48.600 0.700 ;
        RECT 49.000 0.300 49.400 0.700 ;
      LAYER metal4 ;
        RECT 48.000 120.300 49.600 120.700 ;
        RECT 48.000 100.300 49.600 100.700 ;
        RECT 48.000 80.300 49.600 80.700 ;
        RECT 48.000 60.300 49.600 60.700 ;
        RECT 48.000 40.300 49.600 40.700 ;
        RECT 48.000 20.300 49.600 20.700 ;
        RECT 48.000 0.300 49.600 0.700 ;
      LAYER via4 ;
        RECT 48.200 120.300 48.600 120.700 ;
        RECT 48.900 120.300 49.300 120.700 ;
        RECT 48.200 100.300 48.600 100.700 ;
        RECT 48.900 100.300 49.300 100.700 ;
        RECT 48.200 80.300 48.600 80.700 ;
        RECT 48.900 80.300 49.300 80.700 ;
        RECT 48.200 60.300 48.600 60.700 ;
        RECT 48.900 60.300 49.300 60.700 ;
        RECT 48.200 40.300 48.600 40.700 ;
        RECT 48.900 40.300 49.300 40.700 ;
        RECT 48.200 20.300 48.600 20.700 ;
        RECT 48.900 20.300 49.300 20.700 ;
        RECT 48.200 0.300 48.600 0.700 ;
        RECT 48.900 0.300 49.300 0.700 ;
      LAYER metal5 ;
        RECT 48.000 120.200 49.600 120.700 ;
        RECT 48.000 100.200 49.600 100.700 ;
        RECT 48.000 80.200 49.600 80.700 ;
        RECT 48.000 60.200 49.600 60.700 ;
        RECT 48.000 40.200 49.600 40.700 ;
        RECT 48.000 20.200 49.600 20.700 ;
        RECT 48.000 0.200 49.600 0.700 ;
      LAYER via5 ;
        RECT 49.000 120.200 49.500 120.700 ;
        RECT 49.000 100.200 49.500 100.700 ;
        RECT 49.000 80.200 49.500 80.700 ;
        RECT 49.000 60.200 49.500 60.700 ;
        RECT 49.000 40.200 49.500 40.700 ;
        RECT 49.000 20.200 49.500 20.700 ;
        RECT 49.000 0.200 49.500 0.700 ;
      LAYER metal6 ;
        RECT 48.000 -3.000 49.600 133.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.200 130.200 151.000 130.800 ;
        RECT 3.000 126.900 3.400 130.200 ;
        RECT 4.100 127.900 4.500 130.200 ;
        RECT 6.200 128.900 6.600 130.200 ;
        RECT 7.000 128.900 7.400 130.200 ;
        RECT 9.100 127.900 9.500 130.200 ;
        RECT 10.200 126.900 10.600 130.200 ;
        RECT 14.200 128.300 14.600 130.200 ;
        RECT 19.000 126.900 19.400 130.200 ;
        RECT 20.600 128.300 21.000 130.200 ;
        RECT 23.000 126.900 23.400 130.200 ;
        RECT 26.200 127.900 26.600 130.200 ;
        RECT 29.200 127.900 29.600 130.200 ;
        RECT 30.200 128.900 30.600 130.200 ;
        RECT 31.800 128.900 32.200 130.200 ;
        RECT 33.400 128.900 33.800 130.200 ;
        RECT 35.000 129.100 35.400 130.200 ;
        RECT 41.400 126.900 41.800 130.200 ;
        RECT 43.000 128.300 43.400 130.200 ;
        RECT 45.700 127.900 46.100 130.200 ;
        RECT 47.800 128.900 48.200 130.200 ;
        RECT 50.200 126.900 50.600 130.200 ;
        RECT 55.800 126.900 56.200 130.200 ;
        RECT 59.800 129.100 60.200 130.200 ;
        RECT 61.400 128.900 61.800 130.200 ;
        RECT 63.800 128.300 64.200 130.200 ;
        RECT 66.200 128.900 66.600 130.200 ;
        RECT 67.800 126.900 68.200 130.200 ;
        RECT 71.800 128.900 72.200 130.200 ;
        RECT 75.000 126.900 75.400 130.200 ;
        RECT 75.800 127.900 76.200 130.200 ;
        RECT 77.400 127.900 77.800 130.200 ;
        RECT 79.000 127.900 79.400 130.200 ;
        RECT 82.200 126.900 82.600 130.200 ;
        RECT 84.600 127.900 85.000 130.200 ;
        RECT 89.400 128.900 89.800 130.200 ;
        RECT 91.000 128.900 91.400 130.200 ;
        RECT 96.600 127.900 97.000 130.200 ;
        RECT 99.800 128.900 100.200 130.200 ;
        RECT 103.800 127.900 104.200 130.200 ;
        RECT 108.600 128.900 109.000 130.200 ;
        RECT 110.200 128.900 110.600 130.200 ;
        RECT 115.800 127.900 116.200 130.200 ;
        RECT 119.000 128.900 119.400 130.200 ;
        RECT 120.600 128.900 121.000 130.200 ;
        RECT 123.000 127.900 123.400 130.200 ;
        RECT 127.800 128.900 128.200 130.200 ;
        RECT 129.400 128.900 129.800 130.200 ;
        RECT 135.000 127.900 135.400 130.200 ;
        RECT 138.200 128.900 138.600 130.200 ;
        RECT 139.800 127.900 140.200 130.200 ;
        RECT 142.200 127.900 142.600 130.200 ;
        RECT 144.600 127.900 145.000 130.200 ;
        RECT 146.200 127.900 146.600 130.200 ;
        RECT 149.400 127.900 149.800 130.200 ;
        RECT 3.000 110.800 3.400 114.100 ;
        RECT 6.200 110.800 6.600 114.100 ;
        RECT 7.000 110.800 7.400 112.100 ;
        RECT 8.600 110.800 9.000 112.100 ;
        RECT 11.800 110.800 12.200 114.100 ;
        RECT 14.200 110.800 14.600 113.100 ;
        RECT 15.000 110.800 15.400 114.100 ;
        RECT 19.800 110.800 20.200 112.700 ;
        RECT 22.200 110.800 22.600 113.100 ;
        RECT 23.300 110.800 23.700 113.100 ;
        RECT 25.400 110.800 25.800 112.100 ;
        RECT 27.000 110.800 27.400 112.700 ;
        RECT 29.700 110.800 30.100 113.100 ;
        RECT 31.800 110.800 32.200 112.100 ;
        RECT 35.000 110.800 35.400 114.100 ;
        RECT 35.800 110.800 36.200 114.100 ;
        RECT 40.600 110.800 41.000 112.700 ;
        RECT 42.200 110.800 42.600 114.100 ;
        RECT 45.400 110.800 45.800 112.100 ;
        RECT 47.500 110.800 47.900 113.100 ;
        RECT 51.000 110.800 51.400 112.100 ;
        RECT 51.800 110.800 52.200 113.100 ;
        RECT 54.200 110.800 54.600 112.100 ;
        RECT 55.800 110.800 56.200 112.100 ;
        RECT 56.600 110.800 57.000 112.100 ;
        RECT 58.200 110.800 58.600 112.900 ;
        RECT 59.800 110.800 60.200 112.100 ;
        RECT 61.900 110.800 62.300 113.100 ;
        RECT 63.800 110.800 64.200 113.100 ;
        RECT 64.600 110.800 65.000 112.100 ;
        RECT 66.700 110.800 67.100 113.100 ;
        RECT 67.800 110.800 68.200 114.100 ;
        RECT 71.800 110.800 72.200 112.700 ;
        RECT 76.600 110.800 77.000 114.100 ;
        RECT 77.400 110.800 77.800 112.100 ;
        RECT 79.800 110.800 80.200 112.700 ;
        RECT 83.800 110.800 84.200 113.100 ;
        RECT 88.600 110.800 89.000 112.100 ;
        RECT 90.200 110.800 90.600 112.100 ;
        RECT 95.800 110.800 96.200 113.100 ;
        RECT 99.000 110.800 99.400 112.100 ;
        RECT 101.400 110.800 101.800 112.100 ;
        RECT 103.000 110.800 103.400 112.100 ;
        RECT 103.800 110.800 104.200 113.100 ;
        RECT 105.400 110.800 105.800 113.100 ;
        RECT 108.400 110.800 108.800 113.100 ;
        RECT 111.800 110.800 112.200 114.100 ;
        RECT 113.400 110.800 113.800 112.100 ;
        RECT 114.400 110.800 114.800 113.100 ;
        RECT 117.400 110.800 117.800 113.100 ;
        RECT 118.400 110.800 118.800 113.100 ;
        RECT 121.400 110.800 121.800 113.100 ;
        RECT 123.800 110.800 124.200 113.100 ;
        RECT 128.600 110.800 129.000 112.100 ;
        RECT 130.200 110.800 130.600 112.100 ;
        RECT 135.800 110.800 136.200 113.100 ;
        RECT 139.000 110.800 139.400 112.100 ;
        RECT 140.600 110.800 141.000 112.100 ;
        RECT 142.200 110.800 142.600 113.100 ;
        RECT 144.600 110.800 145.000 113.100 ;
        RECT 147.000 110.800 147.400 113.100 ;
        RECT 0.200 110.200 151.000 110.800 ;
        RECT 2.200 108.300 2.600 110.200 ;
        RECT 3.800 108.900 4.200 110.200 ;
        RECT 5.900 107.900 6.300 110.200 ;
        RECT 9.400 106.900 9.800 110.200 ;
        RECT 10.200 106.900 10.600 110.200 ;
        RECT 13.400 107.900 13.800 110.200 ;
        RECT 15.800 107.900 16.200 110.200 ;
        RECT 17.400 107.900 17.800 110.200 ;
        RECT 22.200 106.900 22.600 110.200 ;
        RECT 25.400 106.900 25.800 110.200 ;
        RECT 26.200 108.900 26.600 110.200 ;
        RECT 28.300 107.900 28.700 110.200 ;
        RECT 29.400 106.900 29.800 110.200 ;
        RECT 32.600 106.900 33.000 110.200 ;
        RECT 35.800 108.900 36.200 110.200 ;
        RECT 37.900 107.900 38.300 110.200 ;
        RECT 39.000 108.900 39.400 110.200 ;
        RECT 41.100 107.900 41.500 110.200 ;
        RECT 42.200 106.900 42.600 110.200 ;
        RECT 45.400 106.900 45.800 110.200 ;
        RECT 50.200 106.900 50.600 110.200 ;
        RECT 55.000 108.300 55.400 110.200 ;
        RECT 58.200 108.300 58.600 110.200 ;
        RECT 60.100 107.900 60.500 110.200 ;
        RECT 62.200 108.900 62.600 110.200 ;
        RECT 63.800 108.300 64.200 110.200 ;
        RECT 67.800 108.300 68.200 110.200 ;
        RECT 71.800 106.900 72.200 110.200 ;
        RECT 72.600 108.900 73.000 110.200 ;
        RECT 74.700 107.900 75.100 110.200 ;
        RECT 75.800 107.900 76.200 110.200 ;
        RECT 79.000 108.900 79.400 110.200 ;
        RECT 79.800 108.900 80.200 110.200 ;
        RECT 81.900 107.900 82.300 110.200 ;
        RECT 83.000 106.900 83.400 110.200 ;
        RECT 86.200 108.900 86.600 110.200 ;
        RECT 88.100 107.900 88.500 110.200 ;
        RECT 90.200 108.900 90.600 110.200 ;
        RECT 91.300 107.900 91.700 110.200 ;
        RECT 93.400 108.900 93.800 110.200 ;
        RECT 94.200 108.900 94.600 110.200 ;
        RECT 95.800 108.900 96.200 110.200 ;
        RECT 96.600 108.900 97.000 110.200 ;
        RECT 98.200 108.900 98.600 110.200 ;
        RECT 99.000 108.900 99.400 110.200 ;
        RECT 100.600 108.900 101.000 110.200 ;
        RECT 104.600 107.900 105.000 110.200 ;
        RECT 109.400 108.900 109.800 110.200 ;
        RECT 111.000 108.900 111.400 110.200 ;
        RECT 116.600 107.900 117.000 110.200 ;
        RECT 119.800 108.900 120.200 110.200 ;
        RECT 122.200 108.300 122.600 110.200 ;
        RECT 125.400 107.900 125.800 110.200 ;
        RECT 130.200 108.900 130.600 110.200 ;
        RECT 131.800 108.900 132.200 110.200 ;
        RECT 137.400 107.900 137.800 110.200 ;
        RECT 140.600 108.900 141.000 110.200 ;
        RECT 141.400 108.900 141.800 110.200 ;
        RECT 143.000 106.900 143.400 110.200 ;
        RECT 146.200 108.900 146.600 110.200 ;
        RECT 147.800 108.900 148.200 110.200 ;
        RECT 3.000 90.800 3.400 94.100 ;
        RECT 3.800 90.800 4.200 93.100 ;
        RECT 7.800 90.800 8.200 94.100 ;
        RECT 8.600 90.800 9.000 93.100 ;
        RECT 11.200 90.800 11.600 93.100 ;
        RECT 14.200 90.800 14.600 93.100 ;
        RECT 17.400 90.800 17.800 94.100 ;
        RECT 18.500 90.800 18.900 93.100 ;
        RECT 20.600 90.800 21.000 92.100 ;
        RECT 22.200 90.800 22.600 92.700 ;
        RECT 24.600 90.800 25.000 92.100 ;
        RECT 26.700 90.800 27.100 93.100 ;
        RECT 30.200 90.800 30.600 94.100 ;
        RECT 33.400 90.800 33.800 94.100 ;
        RECT 34.200 90.800 34.600 92.100 ;
        RECT 36.300 90.800 36.700 93.100 ;
        RECT 37.400 90.800 37.800 94.100 ;
        RECT 41.400 90.800 41.800 93.100 ;
        RECT 42.200 90.800 42.600 94.100 ;
        RECT 45.400 90.800 45.800 94.100 ;
        RECT 50.200 90.800 50.600 94.100 ;
        RECT 53.400 90.800 53.800 94.100 ;
        RECT 56.600 90.800 57.000 92.100 ;
        RECT 58.200 90.800 58.600 92.100 ;
        RECT 61.400 90.800 61.800 94.100 ;
        RECT 62.200 90.800 62.600 92.100 ;
        RECT 64.300 90.800 64.700 93.100 ;
        RECT 65.400 90.800 65.800 92.100 ;
        RECT 67.500 90.800 67.900 93.100 ;
        RECT 68.600 90.800 69.000 94.100 ;
        RECT 71.800 90.800 72.200 92.100 ;
        RECT 73.900 90.800 74.300 93.100 ;
        RECT 75.000 90.800 75.400 92.100 ;
        RECT 76.600 90.800 77.000 92.100 ;
        RECT 78.200 90.800 78.600 92.700 ;
        RECT 83.000 90.800 83.400 92.700 ;
        RECT 85.400 90.800 85.800 92.700 ;
        RECT 88.600 90.800 89.000 93.100 ;
        RECT 91.000 90.800 91.400 92.700 ;
        RECT 92.600 90.800 93.000 92.100 ;
        RECT 94.200 90.800 94.600 92.100 ;
        RECT 97.400 90.800 97.800 94.100 ;
        RECT 99.000 90.800 99.400 92.700 ;
        RECT 103.800 90.800 104.200 92.700 ;
        RECT 107.000 90.800 107.400 92.100 ;
        RECT 107.800 90.800 108.200 92.100 ;
        RECT 109.400 90.800 109.800 92.100 ;
        RECT 110.200 90.800 110.600 92.100 ;
        RECT 111.800 90.800 112.200 92.100 ;
        RECT 114.200 90.800 114.600 93.100 ;
        RECT 115.800 90.800 116.200 92.700 ;
        RECT 118.500 90.800 118.900 93.100 ;
        RECT 120.600 90.800 121.000 92.100 ;
        RECT 121.400 90.800 121.800 92.100 ;
        RECT 123.000 90.800 123.400 92.100 ;
        RECT 125.400 90.800 125.800 93.100 ;
        RECT 130.200 90.800 130.600 92.100 ;
        RECT 131.800 90.800 132.200 92.100 ;
        RECT 137.400 90.800 137.800 93.100 ;
        RECT 140.600 90.800 141.000 92.100 ;
        RECT 142.200 90.800 142.600 93.100 ;
        RECT 143.800 90.800 144.200 92.100 ;
        RECT 145.400 90.800 145.800 92.100 ;
        RECT 147.000 90.800 147.400 93.100 ;
        RECT 148.600 90.800 149.000 92.100 ;
        RECT 0.200 90.200 151.000 90.800 ;
        RECT 0.900 87.900 1.300 90.200 ;
        RECT 3.000 88.900 3.400 90.200 ;
        RECT 5.400 88.300 5.800 90.200 ;
        RECT 9.400 86.900 9.800 90.200 ;
        RECT 10.200 88.900 10.600 90.200 ;
        RECT 12.300 87.900 12.700 90.200 ;
        RECT 15.800 86.900 16.200 90.200 ;
        RECT 16.600 86.900 17.000 90.200 ;
        RECT 20.700 89.900 21.100 90.200 ;
        RECT 20.600 88.200 21.100 89.900 ;
        RECT 23.700 88.200 24.200 90.200 ;
        RECT 27.000 87.900 27.400 90.200 ;
        RECT 29.400 88.300 29.800 90.200 ;
        RECT 32.600 88.300 33.000 90.200 ;
        RECT 36.600 86.900 37.000 90.200 ;
        RECT 37.400 88.900 37.800 90.200 ;
        RECT 39.500 87.900 39.900 90.200 ;
        RECT 42.200 87.900 42.600 90.200 ;
        RECT 44.600 87.900 45.000 90.200 ;
        RECT 47.000 88.300 47.400 90.200 ;
        RECT 50.200 87.900 50.600 90.200 ;
        RECT 53.400 88.300 53.800 90.200 ;
        RECT 56.100 87.900 56.500 90.200 ;
        RECT 58.200 88.900 58.600 90.200 ;
        RECT 60.600 87.900 61.000 90.200 ;
        RECT 63.000 87.900 63.400 90.200 ;
        RECT 65.400 88.300 65.800 90.200 ;
        RECT 68.600 88.300 69.000 90.200 ;
        RECT 71.000 88.300 71.400 90.200 ;
        RECT 75.000 87.900 75.400 90.200 ;
        RECT 76.600 88.200 77.100 90.200 ;
        RECT 79.700 89.900 80.100 90.200 ;
        RECT 79.700 88.200 80.200 89.900 ;
        RECT 82.700 88.000 83.100 90.200 ;
        RECT 85.400 87.900 85.800 90.200 ;
        RECT 86.200 87.900 86.600 90.200 ;
        RECT 87.800 87.900 88.200 90.200 ;
        RECT 89.400 88.300 89.800 90.200 ;
        RECT 91.800 88.900 92.200 90.200 ;
        RECT 93.900 87.900 94.300 90.200 ;
        RECT 95.000 88.900 95.400 90.200 ;
        RECT 96.600 88.900 97.000 90.200 ;
        RECT 97.400 88.900 97.800 90.200 ;
        RECT 101.400 88.200 101.900 90.200 ;
        RECT 104.500 89.900 104.900 90.200 ;
        RECT 104.500 88.200 105.000 89.900 ;
        RECT 107.800 87.900 108.200 90.200 ;
        RECT 108.600 87.900 109.000 90.200 ;
        RECT 110.200 87.900 110.600 90.200 ;
        RECT 111.300 87.900 111.700 90.200 ;
        RECT 113.400 88.900 113.800 90.200 ;
        RECT 115.800 88.300 116.200 90.200 ;
        RECT 117.400 88.900 117.800 90.200 ;
        RECT 119.000 88.900 119.400 90.200 ;
        RECT 119.800 88.900 120.200 90.200 ;
        RECT 121.400 88.100 121.800 90.200 ;
        RECT 123.300 87.900 123.700 90.200 ;
        RECT 125.400 88.900 125.800 90.200 ;
        RECT 127.000 88.300 127.400 90.200 ;
        RECT 130.200 88.300 130.600 90.200 ;
        RECT 133.500 89.900 133.900 90.200 ;
        RECT 133.400 88.200 133.900 89.900 ;
        RECT 136.500 88.200 137.000 90.200 ;
        RECT 138.500 87.900 138.900 90.200 ;
        RECT 140.600 88.900 141.000 90.200 ;
        RECT 143.000 88.300 143.400 90.200 ;
        RECT 145.400 88.900 145.800 90.200 ;
        RECT 147.000 87.900 147.400 90.200 ;
        RECT 150.200 87.900 150.600 90.200 ;
        RECT 3.000 70.800 3.400 74.100 ;
        RECT 5.400 70.800 5.800 72.700 ;
        RECT 9.400 70.800 9.800 74.100 ;
        RECT 10.200 70.800 10.600 72.100 ;
        RECT 12.300 70.800 12.700 73.100 ;
        RECT 13.400 70.800 13.800 74.100 ;
        RECT 18.200 70.800 18.600 73.100 ;
        RECT 19.800 70.800 20.200 72.700 ;
        RECT 23.000 70.800 23.400 72.700 ;
        RECT 27.000 70.800 27.400 73.100 ;
        RECT 27.800 70.800 28.200 72.100 ;
        RECT 31.000 70.800 31.400 72.700 ;
        RECT 33.400 70.800 33.800 72.700 ;
        RECT 37.400 70.800 37.800 73.100 ;
        RECT 38.200 70.800 38.600 72.100 ;
        RECT 40.300 70.800 40.700 73.100 ;
        RECT 43.800 70.800 44.200 74.100 ;
        RECT 44.600 70.800 45.000 72.100 ;
        RECT 46.700 70.800 47.100 73.100 ;
        RECT 49.400 70.800 49.800 74.100 ;
        RECT 53.400 70.800 53.800 72.100 ;
        RECT 54.200 70.800 54.600 74.100 ;
        RECT 57.400 70.800 57.800 74.100 ;
        RECT 60.600 70.800 61.000 72.100 ;
        RECT 62.200 70.800 62.600 72.100 ;
        RECT 64.600 70.800 65.000 72.700 ;
        RECT 67.000 70.800 67.400 72.700 ;
        RECT 69.400 70.800 69.800 72.100 ;
        RECT 71.000 70.800 71.400 72.100 ;
        RECT 72.600 70.800 73.000 72.700 ;
        RECT 75.000 70.800 75.400 73.100 ;
        RECT 76.600 70.800 77.000 73.100 ;
        RECT 79.000 70.800 79.400 73.100 ;
        RECT 80.600 70.800 81.000 73.100 ;
        RECT 81.400 70.800 81.800 73.100 ;
        RECT 84.600 70.800 85.000 72.700 ;
        RECT 87.000 70.800 87.400 72.100 ;
        RECT 88.600 70.800 89.000 72.100 ;
        RECT 90.200 70.800 90.600 72.700 ;
        RECT 92.600 70.800 93.000 73.100 ;
        RECT 96.300 70.800 96.700 73.000 ;
        RECT 98.200 70.800 98.600 73.100 ;
        RECT 101.200 70.800 101.600 73.100 ;
        RECT 104.600 70.800 105.000 72.100 ;
        RECT 105.400 70.800 105.800 72.100 ;
        RECT 107.500 70.800 107.900 73.100 ;
        RECT 108.900 70.800 109.300 73.100 ;
        RECT 111.000 70.800 111.400 72.100 ;
        RECT 112.900 70.800 113.300 73.000 ;
        RECT 115.000 70.800 115.400 72.100 ;
        RECT 116.600 70.800 117.000 72.100 ;
        RECT 119.000 70.800 119.400 72.700 ;
        RECT 122.200 70.800 122.600 73.100 ;
        RECT 123.000 70.800 123.400 72.100 ;
        RECT 125.100 70.800 125.500 73.100 ;
        RECT 127.500 70.800 127.900 73.000 ;
        RECT 129.400 70.800 129.800 72.100 ;
        RECT 131.000 70.800 131.400 72.100 ;
        RECT 131.800 70.800 132.200 73.100 ;
        RECT 134.200 70.800 134.600 72.700 ;
        RECT 137.400 70.800 137.800 72.700 ;
        RECT 141.400 70.800 141.800 72.700 ;
        RECT 143.000 70.800 143.400 72.100 ;
        RECT 144.600 70.800 145.000 72.900 ;
        RECT 147.000 70.800 147.400 73.100 ;
        RECT 147.800 70.800 148.200 73.100 ;
        RECT 0.200 70.200 151.000 70.800 ;
        RECT 0.900 67.900 1.300 70.200 ;
        RECT 3.000 68.900 3.400 70.200 ;
        RECT 3.800 68.900 4.200 70.200 ;
        RECT 5.400 68.900 5.800 70.200 ;
        RECT 6.200 68.900 6.600 70.200 ;
        RECT 8.300 67.900 8.700 70.200 ;
        RECT 9.400 66.900 9.800 70.200 ;
        RECT 15.000 66.900 15.400 70.200 ;
        RECT 15.800 66.900 16.200 70.200 ;
        RECT 20.100 68.000 20.500 70.200 ;
        RECT 22.200 68.900 22.600 70.200 ;
        RECT 23.800 68.900 24.200 70.200 ;
        RECT 27.000 68.300 27.400 70.200 ;
        RECT 30.200 67.900 30.600 70.200 ;
        RECT 31.000 68.900 31.400 70.200 ;
        RECT 33.100 67.900 33.500 70.200 ;
        RECT 35.800 67.900 36.200 70.200 ;
        RECT 38.200 67.900 38.600 70.200 ;
        RECT 40.600 68.300 41.000 70.200 ;
        RECT 43.000 68.300 43.400 70.200 ;
        RECT 47.000 68.300 47.400 70.200 ;
        RECT 51.000 68.300 51.400 70.200 ;
        RECT 55.000 67.900 55.400 70.200 ;
        RECT 56.600 68.300 57.000 70.200 ;
        RECT 59.800 67.900 60.200 70.200 ;
        RECT 62.800 67.900 63.200 70.200 ;
        RECT 63.800 68.900 64.200 70.200 ;
        RECT 65.900 67.900 66.300 70.200 ;
        RECT 67.300 67.900 67.700 70.200 ;
        RECT 69.400 68.900 69.800 70.200 ;
        RECT 70.200 67.900 70.600 70.200 ;
        RECT 74.200 67.900 74.600 70.200 ;
        RECT 75.800 68.300 76.200 70.200 ;
        RECT 79.000 67.700 79.400 70.200 ;
        RECT 81.600 67.500 82.000 70.200 ;
        RECT 83.000 67.900 83.400 70.200 ;
        RECT 85.400 67.900 85.800 70.200 ;
        RECT 87.800 68.900 88.200 70.200 ;
        RECT 89.400 68.900 89.800 70.200 ;
        RECT 90.200 68.900 90.600 70.200 ;
        RECT 92.600 68.300 93.000 70.200 ;
        RECT 95.000 68.900 95.400 70.200 ;
        RECT 96.600 68.900 97.000 70.200 ;
        RECT 97.400 68.900 97.800 70.200 ;
        RECT 99.000 68.900 99.400 70.200 ;
        RECT 102.200 68.300 102.600 70.200 ;
        RECT 104.600 67.900 105.000 70.200 ;
        RECT 108.600 68.300 109.000 70.200 ;
        RECT 111.800 68.300 112.200 70.200 ;
        RECT 113.400 68.900 113.800 70.200 ;
        RECT 115.000 68.900 115.400 70.200 ;
        RECT 116.600 68.300 117.000 70.200 ;
        RECT 119.000 68.900 119.400 70.200 ;
        RECT 120.600 68.900 121.000 70.200 ;
        RECT 121.400 67.900 121.800 70.200 ;
        RECT 125.400 68.300 125.800 70.200 ;
        RECT 127.000 68.900 127.400 70.200 ;
        RECT 128.600 67.900 129.000 70.200 ;
        RECT 131.000 68.900 131.400 70.200 ;
        RECT 132.800 67.900 133.200 70.200 ;
        RECT 135.800 67.900 136.200 70.200 ;
        RECT 136.600 67.900 137.000 70.200 ;
        RECT 139.600 67.900 140.000 70.200 ;
        RECT 140.600 66.900 141.000 70.200 ;
        RECT 144.600 68.100 145.000 70.200 ;
        RECT 146.200 68.900 146.600 70.200 ;
        RECT 147.000 68.900 147.400 70.200 ;
        RECT 149.100 67.900 149.500 70.200 ;
        RECT 0.600 50.800 1.000 52.100 ;
        RECT 2.200 50.800 2.600 54.100 ;
        RECT 6.200 50.800 6.600 52.900 ;
        RECT 7.800 50.800 8.200 52.100 ;
        RECT 10.200 50.800 10.600 52.700 ;
        RECT 13.400 50.800 13.800 52.700 ;
        RECT 15.300 50.800 15.700 53.100 ;
        RECT 17.400 50.800 17.800 52.100 ;
        RECT 18.200 50.800 18.600 54.100 ;
        RECT 23.800 50.800 24.200 54.100 ;
        RECT 27.000 50.800 27.400 54.100 ;
        RECT 27.800 50.800 28.200 52.100 ;
        RECT 29.900 50.800 30.300 53.100 ;
        RECT 31.000 50.800 31.400 54.100 ;
        RECT 34.200 50.800 34.600 54.100 ;
        RECT 38.200 50.800 38.600 52.700 ;
        RECT 41.400 50.800 41.800 53.100 ;
        RECT 44.400 50.800 44.800 53.100 ;
        RECT 45.400 50.800 45.800 52.100 ;
        RECT 47.500 50.800 47.900 53.100 ;
        RECT 51.000 50.800 51.400 53.100 ;
        RECT 51.800 50.800 52.200 52.100 ;
        RECT 53.900 50.800 54.300 53.100 ;
        RECT 55.000 50.800 55.400 52.100 ;
        RECT 56.600 50.800 57.000 52.100 ;
        RECT 57.400 50.800 57.800 52.100 ;
        RECT 59.500 50.800 59.900 53.100 ;
        RECT 60.600 50.800 61.000 53.100 ;
        RECT 63.000 50.800 63.400 53.100 ;
        RECT 64.600 50.800 65.000 53.100 ;
        RECT 66.200 50.800 66.600 53.100 ;
        RECT 67.000 50.800 67.400 52.100 ;
        RECT 68.600 50.800 69.000 52.100 ;
        RECT 69.400 50.800 69.800 52.100 ;
        RECT 71.000 50.800 71.400 52.100 ;
        RECT 72.600 50.800 73.000 52.100 ;
        RECT 73.400 50.800 73.800 52.100 ;
        RECT 75.000 50.800 75.400 52.100 ;
        RECT 76.600 50.800 77.000 53.100 ;
        RECT 79.000 50.800 79.400 52.700 ;
        RECT 80.600 50.800 81.000 53.100 ;
        RECT 83.000 50.800 83.400 52.100 ;
        RECT 84.600 50.800 85.000 52.100 ;
        RECT 86.200 50.800 86.600 52.700 ;
        RECT 88.600 50.800 89.000 52.100 ;
        RECT 91.000 50.800 91.400 52.700 ;
        RECT 94.200 50.800 94.600 52.700 ;
        RECT 96.600 50.800 97.000 52.100 ;
        RECT 98.200 50.800 98.600 52.100 ;
        RECT 101.400 50.800 101.800 52.700 ;
        RECT 103.800 50.800 104.200 52.100 ;
        RECT 105.400 50.800 105.800 52.100 ;
        RECT 107.000 50.800 107.400 52.100 ;
        RECT 107.800 50.800 108.200 52.100 ;
        RECT 109.900 50.800 110.300 53.100 ;
        RECT 111.800 50.800 112.200 52.700 ;
        RECT 114.200 50.800 114.600 52.100 ;
        RECT 116.600 50.800 117.000 52.700 ;
        RECT 119.000 50.800 119.400 53.100 ;
        RECT 121.400 50.800 121.800 52.100 ;
        RECT 123.000 50.800 123.400 52.100 ;
        RECT 124.100 50.800 124.500 53.100 ;
        RECT 126.200 50.800 126.600 52.100 ;
        RECT 127.800 50.800 128.200 52.700 ;
        RECT 130.200 50.800 130.600 52.100 ;
        RECT 132.300 50.800 132.700 53.100 ;
        RECT 133.400 50.800 133.800 54.100 ;
        RECT 136.600 50.800 137.000 53.100 ;
        RECT 138.200 50.800 138.600 53.100 ;
        RECT 139.800 50.800 140.200 52.700 ;
        RECT 142.200 50.800 142.600 52.100 ;
        RECT 143.800 50.800 144.200 52.100 ;
        RECT 144.600 50.800 145.000 52.100 ;
        RECT 146.200 50.800 146.600 52.100 ;
        RECT 147.800 50.800 148.200 52.100 ;
        RECT 148.600 50.800 149.000 52.100 ;
        RECT 150.200 50.800 150.600 52.100 ;
        RECT 0.200 50.200 151.000 50.800 ;
        RECT 1.700 48.000 2.100 50.200 ;
        RECT 3.800 47.900 4.200 50.200 ;
        RECT 8.600 46.900 9.000 50.200 ;
        RECT 9.400 47.900 9.800 50.200 ;
        RECT 11.800 48.900 12.200 50.200 ;
        RECT 14.200 48.300 14.600 50.200 ;
        RECT 16.600 48.900 17.000 50.200 ;
        RECT 18.200 48.900 18.600 50.200 ;
        RECT 19.800 48.200 20.300 50.200 ;
        RECT 22.900 49.900 23.300 50.200 ;
        RECT 22.900 48.200 23.400 49.900 ;
        RECT 24.600 48.900 25.000 50.200 ;
        RECT 26.700 47.900 27.100 50.200 ;
        RECT 29.400 48.300 29.800 50.200 ;
        RECT 32.600 48.300 33.000 50.200 ;
        RECT 35.000 48.300 35.400 50.200 ;
        RECT 39.000 48.300 39.400 50.200 ;
        RECT 40.600 48.900 41.000 50.200 ;
        RECT 42.200 48.900 42.600 50.200 ;
        RECT 43.000 48.900 43.400 50.200 ;
        RECT 45.100 47.900 45.500 50.200 ;
        RECT 47.800 47.900 48.200 50.200 ;
        RECT 50.200 48.900 50.600 50.200 ;
        RECT 52.300 47.900 52.700 50.200 ;
        RECT 55.000 47.900 55.400 50.200 ;
        RECT 55.800 47.900 56.200 50.200 ;
        RECT 59.800 48.300 60.200 50.200 ;
        RECT 63.000 47.900 63.400 50.200 ;
        RECT 63.800 47.900 64.200 50.200 ;
        RECT 65.400 47.900 65.800 50.200 ;
        RECT 67.800 47.900 68.200 50.200 ;
        RECT 69.400 47.900 69.800 50.200 ;
        RECT 71.800 47.900 72.200 50.200 ;
        RECT 74.200 47.900 74.600 50.200 ;
        RECT 76.600 48.300 77.000 50.200 ;
        RECT 78.200 48.900 78.600 50.200 ;
        RECT 79.800 48.900 80.200 50.200 ;
        RECT 81.400 48.300 81.800 50.200 ;
        RECT 84.600 48.300 85.000 50.200 ;
        RECT 88.600 48.300 89.000 50.200 ;
        RECT 91.000 48.300 91.400 50.200 ;
        RECT 95.000 47.900 95.400 50.200 ;
        RECT 96.600 48.300 97.000 50.200 ;
        RECT 103.000 48.300 103.400 50.200 ;
        RECT 106.200 48.300 106.600 50.200 ;
        RECT 108.600 48.300 109.000 50.200 ;
        RECT 111.800 48.900 112.200 50.200 ;
        RECT 112.600 48.900 113.000 50.200 ;
        RECT 114.200 48.900 114.600 50.200 ;
        RECT 115.800 48.300 116.200 50.200 ;
        RECT 119.000 48.300 119.400 50.200 ;
        RECT 123.000 47.900 123.400 50.200 ;
        RECT 124.100 47.900 124.500 50.200 ;
        RECT 126.200 48.900 126.600 50.200 ;
        RECT 128.600 48.300 129.000 50.200 ;
        RECT 130.200 46.900 130.600 50.200 ;
        RECT 134.200 47.900 134.600 50.200 ;
        RECT 135.000 48.900 135.400 50.200 ;
        RECT 136.600 48.900 137.000 50.200 ;
        RECT 137.400 47.900 137.800 50.200 ;
        RECT 139.000 47.900 139.400 50.200 ;
        RECT 140.100 47.900 140.500 50.200 ;
        RECT 142.200 48.900 142.600 50.200 ;
        RECT 144.600 47.900 145.000 50.200 ;
        RECT 147.000 48.300 147.400 50.200 ;
        RECT 148.600 48.900 149.000 50.200 ;
        RECT 150.200 48.900 150.600 50.200 ;
        RECT 2.200 30.800 2.600 32.700 ;
        RECT 4.100 30.800 4.500 33.100 ;
        RECT 6.200 30.800 6.600 32.100 ;
        RECT 7.000 30.800 7.400 34.100 ;
        RECT 11.000 30.800 11.400 32.700 ;
        RECT 13.400 30.800 13.800 34.100 ;
        RECT 16.600 30.800 17.000 32.100 ;
        RECT 18.700 30.800 19.100 33.100 ;
        RECT 19.800 30.800 20.200 34.100 ;
        RECT 23.800 31.100 24.300 32.800 ;
        RECT 23.900 30.800 24.300 31.100 ;
        RECT 26.900 30.800 27.400 32.800 ;
        RECT 30.200 30.800 30.600 33.100 ;
        RECT 31.800 30.800 32.200 32.100 ;
        RECT 33.400 30.800 33.800 33.100 ;
        RECT 35.000 30.800 35.400 33.100 ;
        RECT 37.400 30.800 37.800 33.100 ;
        RECT 39.000 30.800 39.400 33.100 ;
        RECT 40.600 30.800 41.000 33.100 ;
        RECT 41.400 30.800 41.800 33.100 ;
        RECT 44.400 30.800 44.800 33.100 ;
        RECT 47.000 30.800 47.400 33.100 ;
        RECT 49.400 30.800 49.800 33.100 ;
        RECT 51.000 30.800 51.400 33.100 ;
        RECT 53.400 30.800 53.800 33.100 ;
        RECT 55.000 30.800 55.400 33.100 ;
        RECT 56.600 30.800 57.000 33.100 ;
        RECT 58.200 30.800 58.600 33.100 ;
        RECT 59.800 30.800 60.200 33.300 ;
        RECT 62.400 30.800 62.800 33.500 ;
        RECT 64.400 30.800 64.800 33.500 ;
        RECT 67.000 30.800 67.400 33.300 ;
        RECT 69.400 30.800 69.800 32.700 ;
        RECT 72.100 30.800 72.500 33.100 ;
        RECT 74.200 30.800 74.600 32.100 ;
        RECT 75.800 30.800 76.200 32.700 ;
        RECT 79.800 30.800 80.200 32.700 ;
        RECT 82.200 30.800 82.600 32.700 ;
        RECT 86.200 30.800 86.600 33.100 ;
        RECT 87.000 30.800 87.400 32.100 ;
        RECT 88.600 30.800 89.000 32.100 ;
        RECT 89.400 30.800 89.800 32.100 ;
        RECT 91.500 30.800 91.900 33.100 ;
        RECT 92.600 30.800 93.000 32.100 ;
        RECT 94.200 30.800 94.600 32.100 ;
        RECT 95.800 30.800 96.200 32.700 ;
        RECT 98.200 30.800 98.600 32.100 ;
        RECT 100.300 30.800 100.700 33.100 ;
        RECT 104.600 30.800 105.000 33.100 ;
        RECT 106.200 30.800 106.600 33.100 ;
        RECT 108.600 30.800 109.000 32.700 ;
        RECT 110.200 30.800 110.600 32.100 ;
        RECT 111.800 30.800 112.200 32.100 ;
        RECT 113.900 30.800 114.300 33.000 ;
        RECT 116.600 30.800 117.000 32.700 ;
        RECT 119.000 30.800 119.400 33.100 ;
        RECT 121.400 30.800 121.800 32.100 ;
        RECT 123.000 30.800 123.400 32.900 ;
        RECT 124.900 30.800 125.300 33.100 ;
        RECT 127.000 30.800 127.400 32.100 ;
        RECT 127.800 30.800 128.200 32.100 ;
        RECT 129.400 30.800 129.800 32.100 ;
        RECT 131.000 30.800 131.400 32.900 ;
        RECT 132.600 30.800 133.000 32.100 ;
        RECT 134.200 30.800 134.600 33.100 ;
        RECT 137.400 30.800 137.800 34.100 ;
        RECT 139.000 30.800 139.400 32.900 ;
        RECT 140.600 30.800 141.000 32.100 ;
        RECT 141.400 30.800 141.800 32.100 ;
        RECT 143.000 30.800 143.400 32.100 ;
        RECT 145.400 30.800 145.800 33.100 ;
        RECT 147.000 30.800 147.400 32.900 ;
        RECT 148.600 30.800 149.000 32.100 ;
        RECT 0.200 30.200 151.000 30.800 ;
        RECT 1.400 28.200 1.900 30.200 ;
        RECT 4.500 29.900 4.900 30.200 ;
        RECT 4.500 28.200 5.000 29.900 ;
        RECT 8.600 26.900 9.000 30.200 ;
        RECT 9.700 27.900 10.100 30.200 ;
        RECT 11.800 28.900 12.200 30.200 ;
        RECT 12.600 28.900 13.000 30.200 ;
        RECT 14.200 28.900 14.600 30.200 ;
        RECT 16.300 27.900 16.700 30.200 ;
        RECT 17.400 26.900 17.800 30.200 ;
        RECT 20.600 27.900 21.000 30.200 ;
        RECT 25.400 26.900 25.800 30.200 ;
        RECT 28.600 26.900 29.000 30.200 ;
        RECT 29.400 27.900 29.800 30.200 ;
        RECT 31.000 27.900 31.400 30.200 ;
        RECT 33.400 27.900 33.800 30.200 ;
        RECT 35.000 27.900 35.400 30.200 ;
        RECT 38.200 28.300 38.600 30.200 ;
        RECT 42.200 26.900 42.600 30.200 ;
        RECT 43.000 26.900 43.400 30.200 ;
        RECT 46.200 27.900 46.600 30.200 ;
        RECT 47.800 27.900 48.200 30.200 ;
        RECT 51.000 27.900 51.400 30.200 ;
        RECT 52.600 27.900 53.000 30.200 ;
        RECT 53.400 27.900 53.800 30.200 ;
        RECT 57.400 28.300 57.800 30.200 ;
        RECT 60.100 28.000 60.500 30.200 ;
        RECT 62.200 28.900 62.600 30.200 ;
        RECT 65.400 27.900 65.800 30.200 ;
        RECT 67.800 28.300 68.200 30.200 ;
        RECT 69.400 27.900 69.800 30.200 ;
        RECT 72.400 27.500 72.800 30.200 ;
        RECT 75.000 27.700 75.400 30.200 ;
        RECT 76.600 28.900 77.000 30.200 ;
        RECT 78.200 28.900 78.600 30.200 ;
        RECT 79.000 28.900 79.400 30.200 ;
        RECT 80.900 27.900 81.300 30.200 ;
        RECT 83.000 28.900 83.400 30.200 ;
        RECT 84.600 28.300 85.000 30.200 ;
        RECT 88.600 28.300 89.000 30.200 ;
        RECT 91.000 28.900 91.400 30.200 ;
        RECT 91.800 28.900 92.200 30.200 ;
        RECT 93.400 28.900 93.800 30.200 ;
        RECT 94.500 27.900 94.900 30.200 ;
        RECT 96.600 28.900 97.000 30.200 ;
        RECT 97.400 27.900 97.800 30.200 ;
        RECT 102.700 28.000 103.100 30.200 ;
        RECT 105.400 28.900 105.800 30.200 ;
        RECT 107.800 28.300 108.200 30.200 ;
        RECT 109.700 27.900 110.100 30.200 ;
        RECT 111.800 28.900 112.200 30.200 ;
        RECT 112.900 27.900 113.300 30.200 ;
        RECT 115.000 28.900 115.400 30.200 ;
        RECT 116.100 27.900 116.500 30.200 ;
        RECT 118.200 28.900 118.600 30.200 ;
        RECT 120.600 28.300 121.000 30.200 ;
        RECT 123.800 28.300 124.200 30.200 ;
        RECT 126.700 28.000 127.100 30.200 ;
        RECT 128.600 27.900 129.000 30.200 ;
        RECT 131.000 28.900 131.400 30.200 ;
        RECT 132.600 28.900 133.000 30.200 ;
        RECT 134.200 28.300 134.600 30.200 ;
        RECT 136.900 27.900 137.300 30.200 ;
        RECT 139.000 28.900 139.400 30.200 ;
        RECT 139.800 27.900 140.200 30.200 ;
        RECT 141.400 27.900 141.800 30.200 ;
        RECT 143.000 27.900 143.400 30.200 ;
        RECT 143.800 28.900 144.200 30.200 ;
        RECT 145.400 28.900 145.800 30.200 ;
        RECT 146.200 28.900 146.600 30.200 ;
        RECT 147.800 28.900 148.200 30.200 ;
        RECT 148.600 28.900 149.000 30.200 ;
        RECT 3.000 10.800 3.400 14.100 ;
        RECT 6.200 10.800 6.600 14.100 ;
        RECT 8.600 10.800 9.000 12.700 ;
        RECT 10.200 10.800 10.600 12.100 ;
        RECT 12.300 10.800 12.700 13.100 ;
        RECT 15.000 10.800 15.400 12.700 ;
        RECT 17.400 10.800 17.800 12.700 ;
        RECT 22.200 10.800 22.600 14.100 ;
        RECT 23.000 10.800 23.400 14.100 ;
        RECT 26.200 10.800 26.600 12.100 ;
        RECT 28.300 10.800 28.700 13.100 ;
        RECT 29.400 10.800 29.800 13.100 ;
        RECT 33.100 10.800 33.500 13.000 ;
        RECT 37.400 10.800 37.800 14.100 ;
        RECT 38.200 10.800 38.600 12.100 ;
        RECT 40.300 10.800 40.700 13.100 ;
        RECT 41.400 10.800 41.800 12.100 ;
        RECT 43.800 10.800 44.200 13.100 ;
        RECT 45.400 10.800 45.800 13.100 ;
        RECT 46.200 10.800 46.600 12.100 ;
        RECT 48.300 10.800 48.700 13.100 ;
        RECT 51.300 10.800 51.700 13.100 ;
        RECT 53.400 10.800 53.800 12.100 ;
        RECT 55.000 10.800 55.400 13.100 ;
        RECT 56.600 10.800 57.000 13.100 ;
        RECT 58.000 10.800 58.400 13.500 ;
        RECT 60.600 10.800 61.000 13.300 ;
        RECT 62.200 10.800 62.600 12.100 ;
        RECT 63.800 10.800 64.200 12.100 ;
        RECT 65.400 10.800 65.800 12.100 ;
        RECT 66.200 10.800 66.600 13.100 ;
        RECT 67.800 10.800 68.200 12.100 ;
        RECT 69.400 10.800 69.800 12.100 ;
        RECT 71.000 10.800 71.400 12.700 ;
        RECT 73.400 10.800 73.800 14.100 ;
        RECT 76.600 10.800 77.000 12.100 ;
        RECT 78.200 10.800 78.600 12.100 ;
        RECT 79.800 10.800 80.200 12.100 ;
        RECT 81.400 11.100 81.900 12.800 ;
        RECT 81.500 10.800 81.900 11.100 ;
        RECT 84.500 10.800 85.000 12.800 ;
        RECT 87.800 10.800 88.200 12.700 ;
        RECT 89.400 10.800 89.800 13.100 ;
        RECT 91.300 10.800 91.700 13.100 ;
        RECT 93.400 10.800 93.800 12.100 ;
        RECT 95.800 10.800 96.200 12.700 ;
        RECT 98.500 10.800 98.900 13.000 ;
        RECT 102.200 10.800 102.600 12.100 ;
        RECT 103.800 10.800 104.200 12.100 ;
        RECT 105.400 10.800 105.800 12.700 ;
        RECT 108.600 10.800 109.000 12.700 ;
        RECT 113.400 10.800 113.800 12.700 ;
        RECT 115.000 10.800 115.400 12.100 ;
        RECT 116.600 10.800 117.000 12.100 ;
        RECT 118.500 10.800 118.900 13.000 ;
        RECT 120.600 10.800 121.000 12.100 ;
        RECT 122.200 10.800 122.600 12.100 ;
        RECT 123.800 10.800 124.200 13.100 ;
        RECT 124.600 10.800 125.000 12.100 ;
        RECT 126.200 10.800 126.600 12.100 ;
        RECT 127.000 10.800 127.400 13.100 ;
        RECT 129.400 10.800 129.800 12.700 ;
        RECT 131.800 10.800 132.200 14.100 ;
        RECT 135.000 10.800 135.400 12.100 ;
        RECT 136.600 10.800 137.000 12.100 ;
        RECT 139.800 10.800 140.200 12.700 ;
        RECT 142.200 10.800 142.600 12.100 ;
        RECT 143.800 10.800 144.200 11.900 ;
        RECT 147.800 10.800 148.200 12.100 ;
        RECT 149.400 10.800 149.800 12.100 ;
        RECT 0.200 10.200 151.000 10.800 ;
        RECT 1.500 9.900 1.900 10.200 ;
        RECT 1.400 8.200 1.900 9.900 ;
        RECT 4.500 8.200 5.000 10.200 ;
        RECT 7.100 9.900 7.500 10.200 ;
        RECT 7.000 8.200 7.500 9.900 ;
        RECT 10.100 8.200 10.600 10.200 ;
        RECT 15.000 9.100 15.400 10.200 ;
        RECT 16.600 8.900 17.000 10.200 ;
        RECT 19.000 8.200 19.500 10.200 ;
        RECT 22.100 9.900 22.500 10.200 ;
        RECT 22.100 8.200 22.600 9.900 ;
        RECT 23.800 8.900 24.200 10.200 ;
        RECT 27.000 8.300 27.400 10.200 ;
        RECT 29.500 9.900 29.900 10.200 ;
        RECT 29.400 8.200 29.900 9.900 ;
        RECT 32.500 8.200 33.000 10.200 ;
        RECT 35.000 8.900 35.400 10.200 ;
        RECT 36.600 9.100 37.000 10.200 ;
        RECT 43.800 9.100 44.200 10.200 ;
        RECT 45.400 8.900 45.800 10.200 ;
        RECT 47.800 8.300 48.200 10.200 ;
        RECT 53.400 7.900 53.800 10.200 ;
        RECT 55.000 7.900 55.400 10.200 ;
        RECT 56.600 7.900 57.000 10.200 ;
        RECT 57.400 7.900 57.800 10.200 ;
        RECT 60.600 7.900 61.000 10.200 ;
        RECT 62.200 7.900 62.600 10.200 ;
        RECT 63.000 7.900 63.400 10.200 ;
        RECT 65.400 8.900 65.800 10.200 ;
        RECT 67.000 8.900 67.400 10.200 ;
        RECT 67.800 7.900 68.200 10.200 ;
        RECT 69.400 8.900 69.800 10.200 ;
        RECT 71.000 8.900 71.400 10.200 ;
        RECT 72.600 7.900 73.000 10.200 ;
        RECT 73.400 8.900 73.800 10.200 ;
        RECT 75.000 8.900 75.400 10.200 ;
        RECT 76.600 8.300 77.000 10.200 ;
        RECT 79.800 8.300 80.200 10.200 ;
        RECT 82.200 8.900 82.600 10.200 ;
        RECT 83.800 8.900 84.200 10.200 ;
        RECT 84.600 8.900 85.000 10.200 ;
        RECT 86.200 8.900 86.600 10.200 ;
        RECT 87.800 8.900 88.200 10.200 ;
        RECT 90.200 8.300 90.600 10.200 ;
        RECT 93.400 8.300 93.800 10.200 ;
        RECT 97.400 8.300 97.800 10.200 ;
        RECT 101.400 8.300 101.800 10.200 ;
        RECT 104.600 8.900 105.000 10.200 ;
        RECT 106.200 8.300 106.600 10.200 ;
        RECT 108.600 8.900 109.000 10.200 ;
        RECT 110.200 8.900 110.600 10.200 ;
        RECT 111.000 8.900 111.400 10.200 ;
        RECT 113.400 8.300 113.800 10.200 ;
        RECT 116.600 8.900 117.000 10.200 ;
        RECT 118.200 8.100 118.600 10.200 ;
        RECT 121.400 8.300 121.800 10.200 ;
        RECT 123.000 8.900 123.400 10.200 ;
        RECT 124.600 8.900 125.000 10.200 ;
        RECT 125.400 7.900 125.800 10.200 ;
        RECT 127.800 8.900 128.200 10.200 ;
        RECT 130.200 8.300 130.600 10.200 ;
        RECT 132.600 8.900 133.000 10.200 ;
        RECT 134.200 8.900 134.600 10.200 ;
        RECT 135.000 7.900 135.400 10.200 ;
        RECT 136.600 8.900 137.000 10.200 ;
        RECT 138.200 8.100 138.600 10.200 ;
        RECT 140.100 7.900 140.500 10.200 ;
        RECT 142.200 8.900 142.600 10.200 ;
        RECT 143.300 7.900 143.700 10.200 ;
        RECT 145.400 8.900 145.800 10.200 ;
        RECT 147.000 8.300 147.400 10.200 ;
      LAYER via1 ;
        RECT 100.200 130.300 100.600 130.700 ;
        RECT 100.900 130.300 101.300 130.700 ;
        RECT 100.200 110.300 100.600 110.700 ;
        RECT 100.900 110.300 101.300 110.700 ;
        RECT 100.200 90.300 100.600 90.700 ;
        RECT 100.900 90.300 101.300 90.700 ;
        RECT 100.200 70.300 100.600 70.700 ;
        RECT 100.900 70.300 101.300 70.700 ;
        RECT 100.200 50.300 100.600 50.700 ;
        RECT 100.900 50.300 101.300 50.700 ;
        RECT 100.200 30.300 100.600 30.700 ;
        RECT 100.900 30.300 101.300 30.700 ;
        RECT 100.200 10.300 100.600 10.700 ;
        RECT 100.900 10.300 101.300 10.700 ;
      LAYER metal2 ;
        RECT 100.000 130.300 101.600 130.700 ;
        RECT 100.000 110.300 101.600 110.700 ;
        RECT 100.000 90.300 101.600 90.700 ;
        RECT 100.000 70.300 101.600 70.700 ;
        RECT 100.000 50.300 101.600 50.700 ;
        RECT 100.000 30.300 101.600 30.700 ;
        RECT 100.000 10.300 101.600 10.700 ;
      LAYER via2 ;
        RECT 100.200 130.300 100.600 130.700 ;
        RECT 100.900 130.300 101.300 130.700 ;
        RECT 100.200 110.300 100.600 110.700 ;
        RECT 100.900 110.300 101.300 110.700 ;
        RECT 100.200 90.300 100.600 90.700 ;
        RECT 100.900 90.300 101.300 90.700 ;
        RECT 100.200 70.300 100.600 70.700 ;
        RECT 100.900 70.300 101.300 70.700 ;
        RECT 100.200 50.300 100.600 50.700 ;
        RECT 100.900 50.300 101.300 50.700 ;
        RECT 100.200 30.300 100.600 30.700 ;
        RECT 100.900 30.300 101.300 30.700 ;
        RECT 100.200 10.300 100.600 10.700 ;
        RECT 100.900 10.300 101.300 10.700 ;
      LAYER metal3 ;
        RECT 100.000 130.300 101.600 130.700 ;
        RECT 100.000 110.300 101.600 110.700 ;
        RECT 100.000 90.300 101.600 90.700 ;
        RECT 100.000 70.300 101.600 70.700 ;
        RECT 100.000 50.300 101.600 50.700 ;
        RECT 100.000 30.300 101.600 30.700 ;
        RECT 100.000 10.300 101.600 10.700 ;
      LAYER via3 ;
        RECT 100.200 130.300 100.600 130.700 ;
        RECT 101.000 130.300 101.400 130.700 ;
        RECT 100.200 110.300 100.600 110.700 ;
        RECT 101.000 110.300 101.400 110.700 ;
        RECT 100.200 90.300 100.600 90.700 ;
        RECT 101.000 90.300 101.400 90.700 ;
        RECT 100.200 70.300 100.600 70.700 ;
        RECT 101.000 70.300 101.400 70.700 ;
        RECT 100.200 50.300 100.600 50.700 ;
        RECT 101.000 50.300 101.400 50.700 ;
        RECT 100.200 30.300 100.600 30.700 ;
        RECT 101.000 30.300 101.400 30.700 ;
        RECT 100.200 10.300 100.600 10.700 ;
        RECT 101.000 10.300 101.400 10.700 ;
      LAYER metal4 ;
        RECT 100.000 130.300 101.600 130.700 ;
        RECT 100.000 110.300 101.600 110.700 ;
        RECT 100.000 90.300 101.600 90.700 ;
        RECT 100.000 70.300 101.600 70.700 ;
        RECT 100.000 50.300 101.600 50.700 ;
        RECT 100.000 30.300 101.600 30.700 ;
        RECT 100.000 10.300 101.600 10.700 ;
      LAYER via4 ;
        RECT 100.200 130.300 100.600 130.700 ;
        RECT 100.900 130.300 101.300 130.700 ;
        RECT 100.200 110.300 100.600 110.700 ;
        RECT 100.900 110.300 101.300 110.700 ;
        RECT 100.200 90.300 100.600 90.700 ;
        RECT 100.900 90.300 101.300 90.700 ;
        RECT 100.200 70.300 100.600 70.700 ;
        RECT 100.900 70.300 101.300 70.700 ;
        RECT 100.200 50.300 100.600 50.700 ;
        RECT 100.900 50.300 101.300 50.700 ;
        RECT 100.200 30.300 100.600 30.700 ;
        RECT 100.900 30.300 101.300 30.700 ;
        RECT 100.200 10.300 100.600 10.700 ;
        RECT 100.900 10.300 101.300 10.700 ;
      LAYER metal5 ;
        RECT 100.000 130.200 101.600 130.700 ;
        RECT 100.000 110.200 101.600 110.700 ;
        RECT 100.000 90.200 101.600 90.700 ;
        RECT 100.000 70.200 101.600 70.700 ;
        RECT 100.000 50.200 101.600 50.700 ;
        RECT 100.000 30.200 101.600 30.700 ;
        RECT 100.000 10.200 101.600 10.700 ;
      LAYER via5 ;
        RECT 101.000 130.200 101.500 130.700 ;
        RECT 101.000 110.200 101.500 110.700 ;
        RECT 101.000 90.200 101.500 90.700 ;
        RECT 101.000 70.200 101.500 70.700 ;
        RECT 101.000 50.200 101.500 50.700 ;
        RECT 101.000 30.200 101.500 30.700 ;
        RECT 101.000 10.200 101.500 10.700 ;
      LAYER metal6 ;
        RECT 100.000 -3.000 101.600 133.000 ;
    END
  END gnd
  PIN a[0]
    PORT
      LAYER metal1 ;
        RECT 60.600 86.800 61.000 87.600 ;
        RECT 75.000 86.800 75.400 87.600 ;
        RECT 86.200 86.800 86.600 87.600 ;
        RECT 55.000 66.800 55.400 67.600 ;
        RECT 85.400 66.800 85.800 67.600 ;
        RECT 84.600 52.400 85.000 53.200 ;
        RECT 57.400 6.800 57.800 7.600 ;
      LAYER via1 ;
        RECT 84.600 52.800 85.000 53.200 ;
      LAYER metal2 ;
        RECT 86.200 87.800 86.600 88.200 ;
        RECT 86.200 87.200 86.500 87.800 ;
        RECT 60.600 86.800 61.000 87.200 ;
        RECT 74.200 87.100 74.600 87.200 ;
        RECT 75.000 87.100 75.400 87.200 ;
        RECT 74.200 86.800 75.400 87.100 ;
        RECT 86.200 86.800 86.600 87.200 ;
        RECT 60.600 81.200 60.900 86.800 ;
        RECT 60.600 80.800 61.000 81.200 ;
        RECT 55.000 67.800 55.400 68.200 ;
        RECT 55.000 67.200 55.300 67.800 ;
        RECT 55.000 66.800 55.400 67.200 ;
        RECT 85.400 66.800 85.800 67.200 ;
        RECT 85.400 66.200 85.700 66.800 ;
        RECT 85.400 65.800 85.800 66.200 ;
        RECT 85.400 55.100 85.700 65.800 ;
        RECT 84.600 54.800 85.700 55.100 ;
        RECT 84.600 53.200 84.900 54.800 ;
        RECT 84.600 52.800 85.000 53.200 ;
        RECT 57.400 28.800 57.800 29.200 ;
        RECT 57.400 7.200 57.700 28.800 ;
        RECT 57.400 6.800 57.800 7.200 ;
        RECT 57.400 -1.800 57.700 6.800 ;
        RECT 57.400 -2.200 57.800 -1.800 ;
      LAYER metal3 ;
        RECT 86.200 87.800 86.600 88.200 ;
        RECT 86.200 87.200 86.500 87.800 ;
        RECT 60.600 87.100 61.000 87.200 ;
        RECT 74.200 87.100 74.600 87.200 ;
        RECT 86.200 87.100 86.600 87.200 ;
        RECT 60.600 86.800 86.600 87.100 ;
        RECT 56.600 81.100 57.000 81.200 ;
        RECT 60.600 81.100 61.000 81.200 ;
        RECT 56.600 80.800 61.000 81.100 ;
        RECT 55.000 67.800 55.400 68.200 ;
        RECT 55.000 67.100 55.300 67.800 ;
        RECT 56.600 67.100 57.000 67.200 ;
        RECT 55.000 66.800 57.000 67.100 ;
        RECT 85.400 66.100 85.800 66.200 ;
        RECT 86.200 66.100 86.600 66.200 ;
        RECT 85.400 65.800 86.600 66.100 ;
        RECT 56.600 29.100 57.000 29.200 ;
        RECT 57.400 29.100 57.800 29.200 ;
        RECT 56.600 28.800 57.800 29.100 ;
      LAYER via3 ;
        RECT 86.200 86.800 86.600 87.200 ;
        RECT 56.600 66.800 57.000 67.200 ;
        RECT 86.200 65.800 86.600 66.200 ;
      LAYER metal4 ;
        RECT 86.200 86.800 86.600 87.200 ;
        RECT 56.600 80.800 57.000 81.200 ;
        RECT 56.600 67.200 56.900 80.800 ;
        RECT 56.600 66.800 57.000 67.200 ;
        RECT 56.600 29.200 56.900 66.800 ;
        RECT 86.200 66.200 86.500 86.800 ;
        RECT 86.200 65.800 86.600 66.200 ;
        RECT 56.600 28.800 57.000 29.200 ;
    END
  END a[0]
  PIN a[1]
    PORT
      LAYER metal1 ;
        RECT 42.200 86.800 42.600 87.600 ;
        RECT 63.000 86.800 63.400 87.600 ;
        RECT 85.400 86.800 85.800 87.600 ;
        RECT 106.200 84.400 106.600 85.200 ;
        RECT 43.800 75.400 44.200 76.200 ;
        RECT 46.600 75.200 47.000 75.400 ;
        RECT 109.000 75.200 109.400 75.400 ;
        RECT 46.600 74.900 47.400 75.200 ;
        RECT 47.000 74.800 47.400 74.900 ;
        RECT 108.600 74.900 109.400 75.200 ;
        RECT 108.600 74.800 109.000 74.900 ;
        RECT 38.200 66.800 38.600 67.600 ;
        RECT 82.200 67.100 82.600 67.200 ;
        RECT 83.000 67.100 83.400 67.600 ;
        RECT 82.200 66.800 83.400 67.100 ;
        RECT 82.200 55.800 82.600 57.200 ;
        RECT 138.200 54.100 138.600 54.200 ;
        RECT 139.000 54.100 139.400 54.200 ;
        RECT 138.200 53.800 139.800 54.100 ;
        RECT 139.400 53.600 139.800 53.800 ;
      LAYER via1 ;
        RECT 106.200 84.800 106.600 85.200 ;
        RECT 43.800 75.800 44.200 76.200 ;
        RECT 82.200 56.800 82.600 57.200 ;
      LAYER metal2 ;
        RECT 42.200 86.800 42.600 87.200 ;
        RECT 63.000 86.800 63.400 87.200 ;
        RECT 85.400 86.800 85.800 87.200 ;
        RECT 42.200 86.200 42.500 86.800 ;
        RECT 63.000 86.200 63.300 86.800 ;
        RECT 42.200 85.800 42.600 86.200 ;
        RECT 47.000 85.800 47.400 86.200 ;
        RECT 63.000 85.800 63.400 86.200 ;
        RECT 43.800 75.800 44.200 76.200 ;
        RECT 43.800 75.200 44.100 75.800 ;
        RECT 47.000 75.200 47.300 85.800 ;
        RECT 63.000 83.200 63.300 85.800 ;
        RECT 85.400 84.200 85.700 86.800 ;
        RECT 106.200 84.800 106.600 85.200 ;
        RECT 106.200 84.200 106.500 84.800 ;
        RECT 85.400 83.800 85.800 84.200 ;
        RECT 106.200 83.800 106.600 84.200 ;
        RECT 63.000 82.800 63.400 83.200 ;
        RECT 106.200 75.200 106.500 83.800 ;
        RECT 108.600 75.800 109.000 76.200 ;
        RECT 108.600 75.200 108.900 75.800 ;
        RECT 43.800 74.800 44.200 75.200 ;
        RECT 47.000 74.800 47.400 75.200 ;
        RECT 106.200 74.800 106.600 75.200 ;
        RECT 108.600 74.800 109.000 75.200 ;
        RECT 138.200 74.800 138.600 75.200 ;
        RECT 47.000 67.200 47.300 74.800 ;
        RECT 82.200 68.800 82.600 69.200 ;
        RECT 82.200 67.200 82.500 68.800 ;
        RECT 38.200 67.100 38.600 67.200 ;
        RECT 39.000 67.100 39.400 67.200 ;
        RECT 38.200 66.800 39.400 67.100 ;
        RECT 47.000 66.800 47.400 67.200 ;
        RECT 82.200 66.800 82.600 67.200 ;
        RECT 82.200 57.200 82.500 66.800 ;
        RECT 82.200 56.800 82.600 57.200 ;
        RECT 138.200 56.200 138.500 74.800 ;
        RECT 138.200 55.800 138.600 56.200 ;
        RECT 138.200 54.200 138.500 55.800 ;
        RECT 138.200 53.800 138.600 54.200 ;
      LAYER via2 ;
        RECT 39.000 66.800 39.400 67.200 ;
      LAYER metal3 ;
        RECT 42.200 86.100 42.600 86.200 ;
        RECT 47.000 86.100 47.400 86.200 ;
        RECT 63.000 86.100 63.400 86.200 ;
        RECT 42.200 85.800 63.400 86.100 ;
        RECT 85.400 84.100 85.800 84.200 ;
        RECT 106.200 84.100 106.600 84.200 ;
        RECT 85.400 83.800 106.600 84.100 ;
        RECT 85.400 83.200 85.700 83.800 ;
        RECT 63.000 83.100 63.400 83.200 ;
        RECT 85.400 83.100 85.800 83.200 ;
        RECT 63.000 82.800 85.800 83.100 ;
        RECT 108.600 75.800 109.000 76.200 ;
        RECT 43.800 75.100 44.200 75.200 ;
        RECT 47.000 75.100 47.400 75.200 ;
        RECT 43.800 74.800 47.400 75.100 ;
        RECT 106.200 75.100 106.600 75.200 ;
        RECT 108.600 75.100 108.900 75.800 ;
        RECT 138.200 75.100 138.600 75.200 ;
        RECT 106.200 74.800 138.600 75.100 ;
        RECT 82.200 69.100 82.600 69.200 ;
        RECT 85.400 69.100 85.800 69.200 ;
        RECT 82.200 68.800 85.800 69.100 ;
        RECT 39.000 67.100 39.400 67.200 ;
        RECT 47.000 67.100 47.400 67.200 ;
        RECT 39.000 66.800 47.400 67.100 ;
        RECT 138.200 56.100 138.600 56.200 ;
        RECT 153.400 56.100 153.800 56.200 ;
        RECT 138.200 55.800 153.800 56.100 ;
      LAYER via3 ;
        RECT 85.400 82.800 85.800 83.200 ;
        RECT 85.400 68.800 85.800 69.200 ;
      LAYER metal4 ;
        RECT 85.400 82.800 85.800 83.200 ;
        RECT 85.400 69.200 85.700 82.800 ;
        RECT 85.400 68.800 85.800 69.200 ;
    END
  END a[1]
  PIN a[2]
    PORT
      LAYER metal1 ;
        RECT 55.800 86.100 56.200 86.200 ;
        RECT 55.800 85.800 56.600 86.100 ;
        RECT 56.200 85.600 56.600 85.800 ;
        RECT 57.400 75.400 57.800 76.200 ;
        RECT 78.200 75.800 78.600 76.600 ;
        RECT 83.000 75.800 83.400 76.600 ;
        RECT 40.200 75.200 40.600 75.400 ;
        RECT 40.200 74.900 41.000 75.200 ;
        RECT 40.600 74.800 41.000 74.900 ;
        RECT 37.400 73.400 37.800 74.200 ;
        RECT 79.000 73.400 79.400 74.200 ;
        RECT 35.800 67.100 36.200 67.600 ;
        RECT 36.600 67.100 37.000 67.200 ;
        RECT 35.800 66.800 37.000 67.100 ;
        RECT 74.200 66.800 74.600 67.600 ;
        RECT 79.000 65.800 79.400 66.600 ;
        RECT 97.400 65.400 97.800 66.200 ;
      LAYER via1 ;
        RECT 57.400 75.800 57.800 76.200 ;
        RECT 37.400 73.800 37.800 74.200 ;
        RECT 79.000 73.800 79.400 74.200 ;
        RECT 36.600 66.800 37.000 67.200 ;
        RECT 97.400 65.800 97.800 66.200 ;
      LAYER metal2 ;
        RECT 55.800 85.800 56.200 86.200 ;
        RECT 55.800 84.200 56.100 85.800 ;
        RECT 55.800 83.800 56.200 84.200 ;
        RECT 57.400 83.800 57.800 84.200 ;
        RECT 57.400 76.200 57.700 83.800 ;
        RECT 37.400 75.800 37.800 76.200 ;
        RECT 40.600 75.800 41.000 76.200 ;
        RECT 57.400 76.100 57.800 76.200 ;
        RECT 58.200 76.100 58.600 76.200 ;
        RECT 57.400 75.800 58.600 76.100 ;
        RECT 78.200 75.800 78.600 76.200 ;
        RECT 82.200 76.100 82.600 76.200 ;
        RECT 83.000 76.100 83.400 76.200 ;
        RECT 82.200 75.800 83.400 76.100 ;
        RECT 37.400 74.200 37.700 75.800 ;
        RECT 40.600 75.200 40.900 75.800 ;
        RECT 40.600 74.800 41.000 75.200 ;
        RECT 37.400 73.800 37.800 74.200 ;
        RECT 78.200 74.100 78.500 75.800 ;
        RECT 83.000 75.200 83.300 75.800 ;
        RECT 83.000 74.800 83.400 75.200 ;
        RECT 97.400 74.800 97.800 75.200 ;
        RECT 79.000 74.100 79.400 74.200 ;
        RECT 78.200 73.800 79.400 74.100 ;
        RECT 36.600 67.100 37.000 67.200 ;
        RECT 37.400 67.100 37.700 73.800 ;
        RECT 79.000 67.200 79.300 73.800 ;
        RECT 36.600 66.800 37.700 67.100 ;
        RECT 73.400 67.100 73.800 67.200 ;
        RECT 74.200 67.100 74.600 67.200 ;
        RECT 73.400 66.800 74.600 67.100 ;
        RECT 79.000 66.800 79.400 67.200 ;
        RECT 79.000 66.200 79.300 66.800 ;
        RECT 97.400 66.200 97.700 74.800 ;
        RECT 79.000 65.800 79.400 66.200 ;
        RECT 97.400 65.800 97.800 66.200 ;
      LAYER via2 ;
        RECT 58.200 75.800 58.600 76.200 ;
      LAYER metal3 ;
        RECT 55.800 84.100 56.200 84.200 ;
        RECT 57.400 84.100 57.800 84.200 ;
        RECT 55.800 83.800 57.800 84.100 ;
        RECT 37.400 76.100 37.800 76.200 ;
        RECT 40.600 76.100 41.000 76.200 ;
        RECT 58.200 76.100 58.600 76.200 ;
        RECT 78.200 76.100 78.600 76.200 ;
        RECT 82.200 76.100 82.600 76.200 ;
        RECT 37.400 75.800 82.600 76.100 ;
        RECT 83.000 75.100 83.400 75.200 ;
        RECT 97.400 75.100 97.800 75.200 ;
        RECT 83.000 74.800 97.800 75.100 ;
        RECT -2.600 67.100 -2.200 67.200 ;
        RECT 0.600 67.100 1.000 67.200 ;
        RECT -2.600 66.800 1.000 67.100 ;
        RECT 35.000 67.100 35.400 67.200 ;
        RECT 36.600 67.100 37.000 67.200 ;
        RECT 35.000 66.800 37.000 67.100 ;
        RECT 73.400 67.100 73.800 67.200 ;
        RECT 79.000 67.100 79.400 67.200 ;
        RECT 73.400 66.800 79.400 67.100 ;
      LAYER via3 ;
        RECT 0.600 66.800 1.000 67.200 ;
      LAYER metal4 ;
        RECT 0.600 67.100 1.000 67.200 ;
        RECT 1.400 67.100 1.800 67.200 ;
        RECT 0.600 66.800 1.800 67.100 ;
        RECT 34.200 67.100 34.600 67.200 ;
        RECT 35.000 67.100 35.400 67.200 ;
        RECT 34.200 66.800 35.400 67.100 ;
      LAYER via4 ;
        RECT 1.400 66.800 1.800 67.200 ;
      LAYER metal5 ;
        RECT 1.400 67.100 1.800 67.200 ;
        RECT 34.200 67.100 34.600 67.200 ;
        RECT 1.400 66.800 34.600 67.100 ;
    END
  END a[2]
  PIN a[3]
    PORT
      LAYER metal1 ;
        RECT 87.800 67.800 88.200 68.600 ;
        RECT 90.200 67.800 90.600 68.600 ;
        RECT 30.200 66.800 30.600 67.600 ;
        RECT 70.200 66.800 70.600 67.600 ;
        RECT 33.400 66.100 33.800 66.200 ;
        RECT 33.000 65.800 33.800 66.100 ;
        RECT 33.000 65.600 33.400 65.800 ;
        RECT 59.800 65.400 60.200 66.200 ;
        RECT 66.200 66.100 66.600 66.200 ;
        RECT 65.800 65.800 66.600 66.100 ;
        RECT 65.800 65.600 66.200 65.800 ;
        RECT 81.400 65.400 81.800 66.200 ;
        RECT 62.200 55.800 62.600 56.600 ;
        RECT 53.400 44.400 53.800 45.200 ;
        RECT 67.000 34.400 67.400 35.200 ;
        RECT 20.600 26.800 21.000 27.600 ;
        RECT 25.400 24.800 25.800 25.600 ;
      LAYER via1 ;
        RECT 33.400 65.800 33.800 66.200 ;
        RECT 59.800 65.800 60.200 66.200 ;
        RECT 66.200 65.800 66.600 66.200 ;
        RECT 81.400 65.800 81.800 66.200 ;
        RECT 53.400 44.800 53.800 45.200 ;
        RECT 67.000 34.800 67.400 35.200 ;
      LAYER metal2 ;
        RECT 87.800 67.800 88.200 68.200 ;
        RECT 90.200 67.800 90.600 68.200 ;
        RECT 30.200 67.100 30.600 67.200 ;
        RECT 31.000 67.100 31.400 67.200 ;
        RECT 30.200 66.800 31.400 67.100 ;
        RECT 33.400 66.800 33.800 67.200 ;
        RECT 70.200 66.800 70.600 67.200 ;
        RECT 33.400 66.200 33.700 66.800 ;
        RECT 33.400 65.800 33.800 66.200 ;
        RECT 59.800 65.800 60.200 66.200 ;
        RECT 66.200 65.800 66.600 66.200 ;
        RECT 33.400 56.200 33.700 65.800 ;
        RECT 59.800 65.200 60.100 65.800 ;
        RECT 66.200 65.200 66.500 65.800 ;
        RECT 70.200 65.200 70.500 66.800 ;
        RECT 87.800 66.200 88.100 67.800 ;
        RECT 90.200 66.200 90.500 67.800 ;
        RECT 81.400 65.800 81.800 66.200 ;
        RECT 87.800 65.800 88.200 66.200 ;
        RECT 90.200 65.800 90.600 66.200 ;
        RECT 59.800 64.800 60.200 65.200 ;
        RECT 66.200 64.800 66.600 65.200 ;
        RECT 70.200 64.800 70.600 65.200 ;
        RECT 59.800 56.200 60.100 64.800 ;
        RECT 81.400 64.200 81.700 65.800 ;
        RECT 87.800 64.200 88.100 65.800 ;
        RECT 81.400 63.800 81.800 64.200 ;
        RECT 87.800 63.800 88.200 64.200 ;
        RECT 33.400 55.800 33.800 56.200 ;
        RECT 59.800 55.800 60.200 56.200 ;
        RECT 61.400 56.100 61.800 56.200 ;
        RECT 62.200 56.100 62.600 56.200 ;
        RECT 61.400 55.800 62.600 56.100 ;
        RECT 20.600 27.800 21.000 28.200 ;
        RECT 20.600 27.200 20.900 27.800 ;
        RECT 20.600 26.800 21.000 27.200 ;
        RECT 20.600 26.200 20.900 26.800 ;
        RECT 33.400 26.200 33.700 55.800 ;
        RECT 62.200 46.200 62.500 55.800 ;
        RECT 53.400 45.800 53.800 46.200 ;
        RECT 62.200 45.800 62.600 46.200 ;
        RECT 67.000 45.800 67.400 46.200 ;
        RECT 53.400 45.200 53.700 45.800 ;
        RECT 53.400 44.800 53.800 45.200 ;
        RECT 67.000 35.200 67.300 45.800 ;
        RECT 67.000 34.800 67.400 35.200 ;
        RECT 20.600 25.800 21.000 26.200 ;
        RECT 25.400 25.800 25.800 26.200 ;
        RECT 33.400 25.800 33.800 26.200 ;
        RECT 25.400 25.200 25.700 25.800 ;
        RECT 25.400 24.800 25.800 25.200 ;
      LAYER via2 ;
        RECT 31.000 66.800 31.400 67.200 ;
      LAYER metal3 ;
        RECT 31.000 67.100 31.400 67.200 ;
        RECT 33.400 67.100 33.800 67.200 ;
        RECT 31.000 66.800 33.800 67.100 ;
        RECT 87.800 66.100 88.200 66.200 ;
        RECT 90.200 66.100 90.600 66.200 ;
        RECT 87.800 65.800 90.600 66.100 ;
        RECT 59.800 65.100 60.200 65.200 ;
        RECT 66.200 65.100 66.600 65.200 ;
        RECT 70.200 65.100 70.600 65.200 ;
        RECT 59.800 64.800 70.600 65.100 ;
        RECT 70.200 64.100 70.500 64.800 ;
        RECT 81.400 64.100 81.800 64.200 ;
        RECT 87.800 64.100 88.200 64.200 ;
        RECT 70.200 63.800 88.200 64.100 ;
        RECT 33.400 56.100 33.800 56.200 ;
        RECT 53.400 56.100 53.800 56.200 ;
        RECT 59.800 56.100 60.200 56.200 ;
        RECT 61.400 56.100 61.800 56.200 ;
        RECT 33.400 55.800 61.800 56.100 ;
        RECT 53.400 46.800 53.800 47.200 ;
        RECT 53.400 46.200 53.700 46.800 ;
        RECT 53.400 45.800 53.800 46.200 ;
        RECT 62.200 46.100 62.600 46.200 ;
        RECT 67.000 46.100 67.400 46.200 ;
        RECT 62.200 45.800 67.400 46.100 ;
        RECT 20.600 28.100 21.000 28.200 ;
        RECT 10.200 27.800 21.000 28.100 ;
        RECT -2.600 27.100 -2.200 27.200 ;
        RECT 10.200 27.100 10.500 27.800 ;
        RECT -2.600 26.800 10.500 27.100 ;
        RECT 20.600 26.100 21.000 26.200 ;
        RECT 25.400 26.100 25.800 26.200 ;
        RECT 33.400 26.100 33.800 26.200 ;
        RECT 20.600 25.800 33.800 26.100 ;
      LAYER via3 ;
        RECT 53.400 55.800 53.800 56.200 ;
      LAYER metal4 ;
        RECT 53.400 55.800 53.800 56.200 ;
        RECT 53.400 47.200 53.700 55.800 ;
        RECT 53.400 46.800 53.800 47.200 ;
    END
  END a[3]
  PIN a[4]
    PORT
      LAYER metal1 ;
        RECT 62.200 66.400 62.600 67.200 ;
        RECT 67.800 66.400 68.200 67.200 ;
        RECT 42.300 54.400 42.700 54.800 ;
        RECT 42.300 54.200 42.600 54.400 ;
        RECT 42.200 53.800 42.600 54.200 ;
        RECT 53.400 53.800 53.800 54.600 ;
        RECT 57.400 44.400 57.800 45.200 ;
        RECT 70.200 44.400 70.600 45.200 ;
        RECT 35.800 35.800 36.200 36.600 ;
        RECT 64.600 34.800 65.000 35.600 ;
        RECT 30.200 33.400 30.600 34.200 ;
        RECT 52.600 26.800 53.000 27.600 ;
        RECT 28.600 24.800 29.000 25.600 ;
        RECT 73.400 14.800 73.800 16.200 ;
        RECT 78.200 12.400 78.600 13.200 ;
      LAYER via1 ;
        RECT 62.200 66.800 62.600 67.200 ;
        RECT 67.800 66.800 68.200 67.200 ;
        RECT 57.400 44.800 57.800 45.200 ;
        RECT 70.200 44.800 70.600 45.200 ;
        RECT 30.200 33.800 30.600 34.200 ;
        RECT 78.200 12.800 78.600 13.200 ;
      LAYER metal2 ;
        RECT 62.200 66.800 62.600 67.200 ;
        RECT 67.000 67.100 67.400 67.200 ;
        RECT 67.800 67.100 68.200 67.200 ;
        RECT 67.000 66.800 68.200 67.100 ;
        RECT 62.200 60.200 62.500 66.800 ;
        RECT 62.200 59.800 62.600 60.200 ;
        RECT 42.200 54.100 42.600 54.200 ;
        RECT 43.000 54.100 43.400 54.200 ;
        RECT 42.200 53.800 43.400 54.100 ;
        RECT 53.400 54.100 53.800 54.200 ;
        RECT 54.200 54.100 54.600 54.200 ;
        RECT 53.400 53.800 54.600 54.100 ;
        RECT 57.400 45.800 57.800 46.200 ;
        RECT 57.400 45.200 57.700 45.800 ;
        RECT 57.400 44.800 57.800 45.200 ;
        RECT 70.200 44.800 70.600 45.200 ;
        RECT 57.400 42.100 57.700 44.800 ;
        RECT 56.600 41.800 57.700 42.100 ;
        RECT 35.800 35.800 36.200 36.200 ;
        RECT 30.200 33.800 30.600 34.200 ;
        RECT 30.200 32.200 30.500 33.800 ;
        RECT 35.800 32.200 36.100 35.800 ;
        RECT 56.600 32.200 56.900 41.800 ;
        RECT 70.200 40.200 70.500 44.800 ;
        RECT 70.200 39.800 70.600 40.200 ;
        RECT 64.600 34.800 65.000 35.200 ;
        RECT 64.600 32.200 64.900 34.800 ;
        RECT 30.200 31.800 30.600 32.200 ;
        RECT 35.800 31.800 36.200 32.200 ;
        RECT 52.600 31.800 53.000 32.200 ;
        RECT 56.600 31.800 57.000 32.200 ;
        RECT 64.600 31.800 65.000 32.200 ;
        RECT 30.200 29.200 30.500 31.800 ;
        RECT 28.600 28.800 29.000 29.200 ;
        RECT 30.200 28.800 30.600 29.200 ;
        RECT 28.600 25.200 28.900 28.800 ;
        RECT 52.600 27.200 52.900 31.800 ;
        RECT 52.600 26.800 53.000 27.200 ;
        RECT 28.600 24.800 29.000 25.200 ;
        RECT 73.400 14.800 73.800 15.200 ;
        RECT 73.400 13.200 73.700 14.800 ;
        RECT 73.400 12.800 73.800 13.200 ;
        RECT 77.400 13.100 77.800 13.200 ;
        RECT 78.200 13.100 78.600 13.200 ;
        RECT 77.400 12.800 78.600 13.100 ;
        RECT 77.400 -0.900 77.700 12.800 ;
        RECT 77.400 -1.200 78.500 -0.900 ;
        RECT 78.200 -1.800 78.500 -1.200 ;
        RECT 78.200 -2.200 78.600 -1.800 ;
      LAYER via2 ;
        RECT 43.000 53.800 43.400 54.200 ;
        RECT 54.200 53.800 54.600 54.200 ;
      LAYER metal3 ;
        RECT 62.200 67.100 62.600 67.200 ;
        RECT 67.000 67.100 67.400 67.200 ;
        RECT 62.200 66.800 67.400 67.100 ;
        RECT 55.800 60.100 56.200 60.200 ;
        RECT 62.200 60.100 62.600 60.200 ;
        RECT 55.800 59.800 62.600 60.100 ;
        RECT 43.000 54.100 43.400 54.200 ;
        RECT 54.200 54.100 54.600 54.200 ;
        RECT 55.800 54.100 56.200 54.200 ;
        RECT 43.000 53.800 56.200 54.100 ;
        RECT 55.800 46.100 56.200 46.200 ;
        RECT 57.400 46.100 57.800 46.200 ;
        RECT 55.800 45.800 57.800 46.100 ;
        RECT 70.200 40.100 70.600 40.200 ;
        RECT 72.600 40.100 73.000 40.200 ;
        RECT 70.200 39.800 73.000 40.100 ;
        RECT 30.200 32.100 30.600 32.200 ;
        RECT 35.800 32.100 36.200 32.200 ;
        RECT 52.600 32.100 53.000 32.200 ;
        RECT 56.600 32.100 57.000 32.200 ;
        RECT 64.600 32.100 65.000 32.200 ;
        RECT 72.600 32.100 73.000 32.200 ;
        RECT 30.200 31.800 73.000 32.100 ;
        RECT 28.600 29.100 29.000 29.200 ;
        RECT 30.200 29.100 30.600 29.200 ;
        RECT 28.600 28.800 30.600 29.100 ;
        RECT 72.600 13.100 73.000 13.200 ;
        RECT 73.400 13.100 73.800 13.200 ;
        RECT 77.400 13.100 77.800 13.200 ;
        RECT 72.600 12.800 77.800 13.100 ;
      LAYER via3 ;
        RECT 55.800 53.800 56.200 54.200 ;
        RECT 72.600 39.800 73.000 40.200 ;
        RECT 72.600 31.800 73.000 32.200 ;
      LAYER metal4 ;
        RECT 55.800 59.800 56.200 60.200 ;
        RECT 55.800 54.200 56.100 59.800 ;
        RECT 55.800 53.800 56.200 54.200 ;
        RECT 55.800 46.200 56.100 53.800 ;
        RECT 55.800 45.800 56.200 46.200 ;
        RECT 72.600 39.800 73.000 40.200 ;
        RECT 72.600 32.200 72.900 39.800 ;
        RECT 72.600 31.800 73.000 32.200 ;
        RECT 72.600 13.200 72.900 31.800 ;
        RECT 72.600 12.800 73.000 13.200 ;
    END
  END a[4]
  PIN a[5]
    PORT
      LAYER metal1 ;
        RECT 43.800 53.800 44.200 54.600 ;
        RECT 59.000 53.800 59.400 54.600 ;
        RECT 51.800 46.400 52.200 47.200 ;
        RECT 46.200 44.400 46.600 45.200 ;
        RECT 61.400 44.400 61.800 45.200 ;
        RECT 42.300 34.400 42.700 34.800 ;
        RECT 42.300 34.200 42.600 34.400 ;
        RECT 42.200 33.800 42.600 34.200 ;
        RECT 60.600 14.400 61.000 15.200 ;
        RECT 66.200 13.400 66.600 14.200 ;
        RECT 65.400 7.800 65.800 8.600 ;
        RECT 51.800 3.800 52.200 5.200 ;
      LAYER via1 ;
        RECT 51.800 46.800 52.200 47.200 ;
        RECT 46.200 44.800 46.600 45.200 ;
        RECT 61.400 44.800 61.800 45.200 ;
        RECT 60.600 14.800 61.000 15.200 ;
        RECT 66.200 13.800 66.600 14.200 ;
      LAYER metal2 ;
        RECT 43.800 53.800 44.200 54.200 ;
        RECT 59.000 53.800 59.400 54.200 ;
        RECT 43.800 51.200 44.100 53.800 ;
        RECT 59.000 51.200 59.300 53.800 ;
        RECT 43.800 50.800 44.200 51.200 ;
        RECT 51.800 50.800 52.200 51.200 ;
        RECT 59.000 50.800 59.400 51.200 ;
        RECT 51.800 47.200 52.100 50.800 ;
        RECT 51.800 46.800 52.200 47.200 ;
        RECT 51.800 45.200 52.100 46.800 ;
        RECT 46.200 44.800 46.600 45.200 ;
        RECT 51.800 44.800 52.200 45.200 ;
        RECT 61.400 44.800 61.800 45.200 ;
        RECT 46.200 34.200 46.500 44.800 ;
        RECT 61.400 44.200 61.700 44.800 ;
        RECT 61.400 43.800 61.800 44.200 ;
        RECT 42.200 34.100 42.600 34.200 ;
        RECT 43.000 34.100 43.400 34.200 ;
        RECT 42.200 33.800 43.400 34.100 ;
        RECT 46.200 33.800 46.600 34.200 ;
        RECT 60.600 14.800 61.000 15.200 ;
        RECT 60.600 8.200 60.900 14.800 ;
        RECT 66.200 13.800 66.600 14.200 ;
        RECT 66.200 12.100 66.500 13.800 ;
        RECT 65.400 11.800 66.500 12.100 ;
        RECT 65.400 8.200 65.700 11.800 ;
        RECT 51.800 7.800 52.200 8.200 ;
        RECT 60.600 7.800 61.000 8.200 ;
        RECT 64.600 8.100 65.000 8.200 ;
        RECT 65.400 8.100 65.800 8.200 ;
        RECT 64.600 7.800 65.800 8.100 ;
        RECT 51.800 4.200 52.100 7.800 ;
        RECT 51.800 3.800 52.200 4.200 ;
        RECT 51.800 -1.800 52.100 3.800 ;
        RECT 51.800 -2.200 52.200 -1.800 ;
      LAYER via2 ;
        RECT 43.000 33.800 43.400 34.200 ;
      LAYER metal3 ;
        RECT 43.800 51.100 44.200 51.200 ;
        RECT 51.800 51.100 52.200 51.200 ;
        RECT 59.000 51.100 59.400 51.200 ;
        RECT 43.800 50.800 59.400 51.100 ;
        RECT 46.200 45.100 46.600 45.200 ;
        RECT 51.800 45.100 52.200 45.200 ;
        RECT 46.200 44.800 52.200 45.100 ;
        RECT 51.800 44.100 52.100 44.800 ;
        RECT 61.400 44.100 61.800 44.200 ;
        RECT 51.800 43.800 61.800 44.100 ;
        RECT 42.200 34.100 42.600 34.200 ;
        RECT 43.000 34.100 43.400 34.200 ;
        RECT 46.200 34.100 46.600 34.200 ;
        RECT 42.200 33.800 46.600 34.100 ;
        RECT 42.200 8.100 42.600 8.200 ;
        RECT 51.800 8.100 52.200 8.200 ;
        RECT 60.600 8.100 61.000 8.200 ;
        RECT 64.600 8.100 65.000 8.200 ;
        RECT 42.200 7.800 65.000 8.100 ;
      LAYER metal4 ;
        RECT 42.200 33.800 42.600 34.200 ;
        RECT 42.200 8.200 42.500 33.800 ;
        RECT 42.200 7.800 42.600 8.200 ;
    END
  END a[5]
  PIN a[6]
    PORT
      LAYER metal1 ;
        RECT 44.600 46.400 45.000 47.200 ;
        RECT 72.600 44.400 73.000 45.200 ;
        RECT 45.400 35.800 45.800 36.600 ;
        RECT 43.800 34.100 44.200 34.600 ;
        RECT 45.400 34.100 45.800 34.200 ;
        RECT 43.800 33.800 45.800 34.100 ;
        RECT 43.800 25.800 44.600 26.200 ;
        RECT 58.200 14.800 58.600 15.600 ;
        RECT 51.800 13.800 52.200 14.600 ;
        RECT 73.400 7.800 73.800 8.600 ;
        RECT 67.800 6.800 68.200 7.600 ;
      LAYER via1 ;
        RECT 44.600 46.800 45.000 47.200 ;
        RECT 72.600 44.800 73.000 45.200 ;
        RECT 45.400 33.800 45.800 34.200 ;
      LAYER metal2 ;
        RECT 44.600 46.800 45.000 47.200 ;
        RECT 44.600 45.100 44.900 46.800 ;
        RECT 44.600 44.800 45.700 45.100 ;
        RECT 45.400 36.200 45.700 44.800 ;
        RECT 72.600 44.800 73.000 45.200 ;
        RECT 45.400 35.800 45.800 36.200 ;
        RECT 45.400 34.200 45.700 35.800 ;
        RECT 43.800 33.800 44.200 34.200 ;
        RECT 45.400 33.800 45.800 34.200 ;
        RECT 43.800 26.200 44.100 33.800 ;
        RECT 72.600 31.200 72.900 44.800 ;
        RECT 72.600 30.800 73.000 31.200 ;
        RECT 43.800 25.800 44.200 26.200 ;
        RECT 43.800 25.200 44.100 25.800 ;
        RECT 43.800 24.800 44.200 25.200 ;
        RECT 51.800 24.800 52.200 25.200 ;
        RECT 51.800 14.200 52.100 24.800 ;
        RECT 58.200 14.800 58.600 15.200 ;
        RECT 51.800 13.800 52.200 14.200 ;
        RECT 51.800 13.200 52.100 13.800 ;
        RECT 58.200 13.200 58.500 14.800 ;
        RECT 51.800 12.800 52.200 13.200 ;
        RECT 58.200 12.800 58.600 13.200 ;
        RECT 67.800 12.800 68.200 13.200 ;
        RECT 67.800 7.200 68.100 12.800 ;
        RECT 73.400 7.800 73.800 8.200 ;
        RECT 73.400 7.200 73.700 7.800 ;
        RECT 67.800 7.100 68.200 7.200 ;
        RECT 68.600 7.100 69.000 7.200 ;
        RECT 67.800 6.800 69.000 7.100 ;
        RECT 73.400 6.800 73.800 7.200 ;
        RECT 68.600 1.200 68.900 6.800 ;
        RECT 68.600 0.800 69.000 1.200 ;
        RECT 70.200 0.800 70.600 1.200 ;
        RECT 70.200 -1.800 70.500 0.800 ;
        RECT 70.200 -2.200 70.600 -1.800 ;
      LAYER via2 ;
        RECT 68.600 6.800 69.000 7.200 ;
      LAYER metal3 ;
        RECT 70.200 31.100 70.600 31.200 ;
        RECT 72.600 31.100 73.000 31.200 ;
        RECT 70.200 30.800 73.000 31.100 ;
        RECT 43.800 25.100 44.200 25.200 ;
        RECT 51.800 25.100 52.200 25.200 ;
        RECT 43.800 24.800 52.200 25.100 ;
        RECT 51.800 13.100 52.200 13.200 ;
        RECT 58.200 13.100 58.600 13.200 ;
        RECT 67.800 13.100 68.200 13.200 ;
        RECT 70.200 13.100 70.600 13.200 ;
        RECT 51.800 12.800 70.600 13.100 ;
        RECT 68.600 7.100 69.000 7.200 ;
        RECT 73.400 7.100 73.800 7.200 ;
        RECT 68.600 6.800 73.800 7.100 ;
        RECT 68.600 1.100 69.000 1.200 ;
        RECT 70.200 1.100 70.600 1.200 ;
        RECT 68.600 0.800 70.600 1.100 ;
      LAYER via3 ;
        RECT 70.200 12.800 70.600 13.200 ;
      LAYER metal4 ;
        RECT 70.200 30.800 70.600 31.200 ;
        RECT 70.200 13.200 70.500 30.800 ;
        RECT 70.200 12.800 70.600 13.200 ;
    END
  END a[6]
  PIN a[7]
    PORT
      LAYER metal1 ;
        RECT 60.400 26.900 60.800 27.000 ;
        RECT 60.400 26.600 60.900 26.900 ;
        RECT 60.600 26.200 60.900 26.600 ;
        RECT 41.000 25.800 41.800 26.200 ;
        RECT 60.600 25.800 61.000 26.200 ;
        RECT 47.800 13.800 48.200 14.600 ;
        RECT 123.000 7.800 123.400 8.600 ;
        RECT 124.600 7.100 125.000 7.200 ;
        RECT 125.400 7.100 125.800 7.600 ;
        RECT 124.600 6.800 125.800 7.100 ;
        RECT 64.600 4.400 65.000 5.200 ;
      LAYER via1 ;
        RECT 41.400 25.800 41.800 26.200 ;
        RECT 64.600 4.800 65.000 5.200 ;
      LAYER metal2 ;
        RECT 41.400 25.800 41.800 26.200 ;
        RECT 60.600 25.800 61.000 26.200 ;
        RECT 41.400 15.200 41.700 25.800 ;
        RECT 60.600 19.200 60.900 25.800 ;
        RECT 47.800 18.800 48.200 19.200 ;
        RECT 60.600 18.800 61.000 19.200 ;
        RECT 47.800 15.200 48.100 18.800 ;
        RECT 41.400 14.800 41.800 15.200 ;
        RECT 47.800 14.800 48.200 15.200 ;
        RECT 47.800 14.200 48.100 14.800 ;
        RECT 47.800 13.800 48.200 14.200 ;
        RECT 123.000 8.100 123.400 8.200 ;
        RECT 123.800 8.100 124.200 8.200 ;
        RECT 123.000 7.800 124.200 8.100 ;
        RECT 124.600 7.800 125.000 8.200 ;
        RECT 124.600 7.200 124.900 7.800 ;
        RECT 124.600 6.800 125.000 7.200 ;
        RECT 63.800 5.100 64.200 5.200 ;
        RECT 64.600 5.100 65.000 5.200 ;
        RECT 63.800 4.800 65.000 5.100 ;
        RECT 66.200 4.800 66.600 5.200 ;
        RECT 66.200 4.200 66.500 4.800 ;
        RECT 124.600 4.200 124.900 6.800 ;
        RECT 66.200 3.800 66.600 4.200 ;
        RECT 124.600 3.800 125.000 4.200 ;
        RECT 66.200 -1.800 66.500 3.800 ;
        RECT 66.200 -2.200 66.600 -1.800 ;
      LAYER via2 ;
        RECT 123.800 7.800 124.200 8.200 ;
      LAYER metal3 ;
        RECT 47.800 19.100 48.200 19.200 ;
        RECT 60.600 19.100 61.000 19.200 ;
        RECT 62.200 19.100 62.600 19.200 ;
        RECT 47.800 18.800 62.600 19.100 ;
        RECT 41.400 15.100 41.800 15.200 ;
        RECT 47.800 15.100 48.200 15.200 ;
        RECT 41.400 14.800 48.200 15.100 ;
        RECT 123.800 8.100 124.200 8.200 ;
        RECT 124.600 8.100 125.000 8.200 ;
        RECT 123.800 7.800 125.000 8.100 ;
        RECT 62.200 5.100 62.600 5.200 ;
        RECT 63.800 5.100 64.200 5.200 ;
        RECT 66.200 5.100 66.600 5.200 ;
        RECT 62.200 4.800 66.600 5.100 ;
        RECT 66.200 4.100 66.600 4.200 ;
        RECT 124.600 4.100 125.000 4.200 ;
        RECT 66.200 3.800 125.000 4.100 ;
      LAYER via3 ;
        RECT 62.200 18.800 62.600 19.200 ;
      LAYER metal4 ;
        RECT 62.200 18.800 62.600 19.200 ;
        RECT 62.200 5.200 62.500 18.800 ;
        RECT 62.200 4.800 62.600 5.200 ;
    END
  END a[7]
  PIN b[0]
    PORT
      LAYER metal1 ;
        RECT 66.100 46.200 66.500 46.600 ;
        RECT 67.100 46.200 67.500 46.600 ;
        RECT 66.100 46.100 66.600 46.200 ;
        RECT 67.000 46.100 67.500 46.200 ;
        RECT 66.100 45.800 67.500 46.100 ;
        RECT 48.500 26.200 48.900 26.600 ;
        RECT 48.500 26.100 49.000 26.200 ;
        RECT 50.200 26.100 50.600 26.200 ;
        RECT 48.500 25.800 50.600 26.100 ;
        RECT 54.200 14.800 54.700 15.200 ;
        RECT 54.300 14.400 54.700 14.800 ;
        RECT 59.900 6.200 60.300 6.600 ;
        RECT 59.800 5.800 60.300 6.200 ;
      LAYER via1 ;
        RECT 66.200 45.800 66.600 46.200 ;
        RECT 50.200 25.800 50.600 26.200 ;
      LAYER metal2 ;
        RECT 66.200 45.800 66.600 46.200 ;
        RECT 66.200 45.200 66.500 45.800 ;
        RECT 66.200 44.800 66.600 45.200 ;
        RECT 50.200 25.800 50.600 26.200 ;
        RECT 50.200 15.200 50.500 25.800 ;
        RECT 50.200 14.800 50.600 15.200 ;
        RECT 54.200 15.100 54.600 15.200 ;
        RECT 55.000 15.100 55.400 15.200 ;
        RECT 54.200 14.800 55.400 15.100 ;
        RECT 59.800 14.800 60.200 15.200 ;
        RECT 59.800 6.200 60.100 14.800 ;
        RECT 59.800 5.800 60.200 6.200 ;
        RECT 59.800 1.200 60.100 5.800 ;
        RECT 59.800 0.800 60.200 1.200 ;
        RECT 63.800 0.800 64.200 1.200 ;
        RECT 63.800 -1.800 64.100 0.800 ;
        RECT 63.800 -2.200 64.200 -1.800 ;
      LAYER via2 ;
        RECT 55.000 14.800 55.400 15.200 ;
      LAYER metal3 ;
        RECT 65.400 45.100 65.800 45.200 ;
        RECT 66.200 45.100 66.600 45.200 ;
        RECT 65.400 44.800 66.600 45.100 ;
        RECT 50.200 15.100 50.600 15.200 ;
        RECT 55.000 15.100 55.400 15.200 ;
        RECT 59.800 15.100 60.200 15.200 ;
        RECT 65.400 15.100 65.800 15.200 ;
        RECT 50.200 14.800 65.800 15.100 ;
        RECT 59.800 1.100 60.200 1.200 ;
        RECT 63.800 1.100 64.200 1.200 ;
        RECT 59.800 0.800 64.200 1.100 ;
      LAYER via3 ;
        RECT 65.400 14.800 65.800 15.200 ;
      LAYER metal4 ;
        RECT 65.400 44.800 65.800 45.200 ;
        RECT 65.400 15.200 65.700 44.800 ;
        RECT 65.400 14.800 65.800 15.200 ;
    END
  END b[0]
  PIN b[1]
    PORT
      LAYER metal1 ;
        RECT 32.600 34.800 33.100 35.200 ;
        RECT 38.200 34.800 38.700 35.200 ;
        RECT 32.700 34.400 33.100 34.800 ;
        RECT 38.300 34.400 38.700 34.800 ;
        RECT 31.700 26.200 32.100 26.600 ;
        RECT 32.700 26.200 33.100 26.600 ;
        RECT 31.700 26.100 32.200 26.200 ;
        RECT 32.600 26.100 33.100 26.200 ;
        RECT 31.700 25.800 33.100 26.100 ;
        RECT 43.000 14.800 43.500 15.200 ;
        RECT 43.100 14.400 43.500 14.800 ;
      LAYER via1 ;
        RECT 32.600 25.800 33.000 26.200 ;
      LAYER metal2 ;
        RECT 32.600 35.800 33.000 36.200 ;
        RECT 38.200 35.800 38.600 36.200 ;
        RECT 32.600 35.200 32.900 35.800 ;
        RECT 38.200 35.200 38.500 35.800 ;
        RECT 32.600 34.800 33.000 35.200 ;
        RECT 38.200 34.800 38.600 35.200 ;
        RECT 32.600 27.800 33.000 28.200 ;
        RECT 32.600 26.200 32.900 27.800 ;
        RECT 32.600 25.800 33.000 26.200 ;
        RECT 32.600 20.200 32.900 25.800 ;
        RECT 32.600 19.800 33.000 20.200 ;
        RECT 43.000 19.800 43.400 20.200 ;
        RECT 43.000 15.200 43.300 19.800 ;
        RECT 43.000 14.800 43.400 15.200 ;
        RECT 43.000 -1.800 43.300 14.800 ;
        RECT 43.000 -2.200 43.400 -1.800 ;
      LAYER metal3 ;
        RECT 32.600 36.100 33.000 36.200 ;
        RECT 38.200 36.100 38.600 36.200 ;
        RECT 32.600 35.800 38.600 36.100 ;
        RECT 32.600 28.800 33.000 29.200 ;
        RECT 32.600 28.200 32.900 28.800 ;
        RECT 32.600 27.800 33.000 28.200 ;
        RECT 32.600 20.100 33.000 20.200 ;
        RECT 43.000 20.100 43.400 20.200 ;
        RECT 32.600 19.800 43.400 20.100 ;
      LAYER metal4 ;
        RECT 32.600 35.800 33.000 36.200 ;
        RECT 32.600 29.200 32.900 35.800 ;
        RECT 32.600 28.800 33.000 29.200 ;
    END
  END b[1]
  PIN b[2]
    PORT
      LAYER metal1 ;
        RECT 51.700 35.100 52.200 35.200 ;
        RECT 52.600 35.100 53.100 35.200 ;
        RECT 51.700 34.800 53.100 35.100 ;
        RECT 55.800 34.800 56.300 35.200 ;
        RECT 51.700 34.400 52.100 34.800 ;
        RECT 52.700 34.400 53.100 34.800 ;
        RECT 55.900 34.400 56.300 34.800 ;
        RECT 54.300 6.200 54.700 6.600 ;
        RECT 54.200 5.800 54.700 6.200 ;
      LAYER via1 ;
        RECT 52.600 34.800 53.000 35.200 ;
      LAYER metal2 ;
        RECT 52.600 34.800 53.000 35.200 ;
        RECT 55.800 34.800 56.200 35.200 ;
        RECT 52.600 34.200 52.900 34.800 ;
        RECT 55.800 34.200 56.100 34.800 ;
        RECT 52.600 33.800 53.000 34.200 ;
        RECT 55.800 33.800 56.200 34.200 ;
        RECT 54.200 5.800 54.600 6.200 ;
        RECT 54.200 -1.800 54.500 5.800 ;
        RECT 54.200 -2.200 54.600 -1.800 ;
      LAYER metal3 ;
        RECT 52.600 34.100 53.000 34.200 ;
        RECT 55.000 34.100 55.400 34.200 ;
        RECT 55.800 34.100 56.200 34.200 ;
        RECT 52.600 33.800 56.200 34.100 ;
        RECT 54.200 6.100 54.600 6.200 ;
        RECT 55.800 6.100 56.200 6.200 ;
        RECT 54.200 5.800 56.200 6.100 ;
      LAYER via3 ;
        RECT 55.000 33.800 55.400 34.200 ;
        RECT 55.800 5.800 56.200 6.200 ;
      LAYER metal4 ;
        RECT 55.000 34.100 55.400 34.200 ;
        RECT 55.000 33.800 56.100 34.100 ;
        RECT 55.800 6.200 56.100 33.800 ;
        RECT 55.800 5.800 56.200 6.200 ;
    END
  END b[2]
  PIN b[3]
    PORT
      LAYER metal1 ;
        RECT 56.600 86.400 57.000 87.200 ;
        RECT 40.600 84.400 41.000 85.200 ;
        RECT 73.400 84.400 73.800 85.200 ;
        RECT 58.200 74.800 59.000 75.200 ;
        RECT 95.000 67.800 95.400 68.600 ;
        RECT 32.600 66.400 33.000 67.200 ;
        RECT 89.400 65.400 89.800 66.200 ;
        RECT 28.600 64.400 29.000 65.200 ;
        RECT 34.200 64.400 34.600 65.200 ;
        RECT 28.600 35.800 29.000 36.600 ;
        RECT 27.400 25.800 28.200 26.200 ;
      LAYER via1 ;
        RECT 56.600 86.800 57.000 87.200 ;
        RECT 40.600 84.800 41.000 85.200 ;
        RECT 73.400 84.800 73.800 85.200 ;
        RECT 32.600 66.800 33.000 67.200 ;
        RECT 89.400 65.800 89.800 66.200 ;
        RECT 28.600 64.800 29.000 65.200 ;
        RECT 34.200 64.800 34.600 65.200 ;
        RECT 27.800 25.800 28.200 26.200 ;
      LAYER metal2 ;
        RECT 56.600 86.800 57.000 87.200 ;
        RECT 40.600 84.800 41.000 85.200 ;
        RECT 40.600 82.200 40.900 84.800 ;
        RECT 56.600 82.200 56.900 86.800 ;
        RECT 73.400 84.800 73.800 85.200 ;
        RECT 73.400 82.200 73.700 84.800 ;
        RECT 32.600 81.800 33.000 82.200 ;
        RECT 40.600 81.800 41.000 82.200 ;
        RECT 56.600 81.800 57.000 82.200 ;
        RECT 73.400 81.800 73.800 82.200 ;
        RECT 32.600 67.200 32.900 81.800 ;
        RECT 56.600 75.200 56.900 81.800 ;
        RECT 56.600 74.800 57.000 75.200 ;
        RECT 57.400 75.100 57.800 75.200 ;
        RECT 58.200 75.100 58.600 75.200 ;
        RECT 57.400 74.800 58.600 75.100 ;
        RECT 89.400 67.800 89.800 68.200 ;
        RECT 94.200 68.100 94.600 68.200 ;
        RECT 95.000 68.100 95.400 68.200 ;
        RECT 94.200 67.800 95.400 68.100 ;
        RECT 32.600 66.800 33.000 67.200 ;
        RECT 32.600 65.200 32.900 66.800 ;
        RECT 89.400 66.200 89.700 67.800 ;
        RECT 89.400 65.800 89.800 66.200 ;
        RECT 28.600 64.800 29.000 65.200 ;
        RECT 32.600 64.800 33.000 65.200 ;
        RECT 34.200 65.100 34.600 65.200 ;
        RECT 35.000 65.100 35.400 65.200 ;
        RECT 34.200 64.800 35.400 65.100 ;
        RECT 28.600 64.200 28.900 64.800 ;
        RECT 28.600 63.800 29.000 64.200 ;
        RECT 28.600 44.800 29.000 45.200 ;
        RECT 28.600 36.200 28.900 44.800 ;
        RECT 28.600 35.800 29.000 36.200 ;
        RECT 28.600 33.100 28.900 35.800 ;
        RECT 27.800 32.800 28.900 33.100 ;
        RECT 27.800 26.200 28.100 32.800 ;
        RECT 27.800 25.800 28.200 26.200 ;
        RECT 27.800 23.200 28.100 25.800 ;
        RECT 27.800 22.800 28.200 23.200 ;
        RECT 27.000 0.800 27.400 1.200 ;
        RECT 27.000 -1.800 27.300 0.800 ;
        RECT 27.000 -2.200 27.400 -1.800 ;
      LAYER via2 ;
        RECT 35.000 64.800 35.400 65.200 ;
      LAYER metal3 ;
        RECT 32.600 82.100 33.000 82.200 ;
        RECT 40.600 82.100 41.000 82.200 ;
        RECT 56.600 82.100 57.000 82.200 ;
        RECT 73.400 82.100 73.800 82.200 ;
        RECT 76.600 82.100 77.000 82.200 ;
        RECT 32.600 81.800 77.000 82.100 ;
        RECT 56.600 75.100 57.000 75.200 ;
        RECT 57.400 75.100 57.800 75.200 ;
        RECT 56.600 74.800 57.800 75.100 ;
        RECT 76.600 68.100 77.000 68.200 ;
        RECT 89.400 68.100 89.800 68.200 ;
        RECT 94.200 68.100 94.600 68.200 ;
        RECT 76.600 67.800 94.600 68.100 ;
        RECT 28.600 65.100 29.000 65.200 ;
        RECT 32.600 65.100 33.000 65.200 ;
        RECT 35.000 65.100 35.400 65.200 ;
        RECT 28.600 64.800 35.400 65.100 ;
        RECT 28.600 64.200 28.900 64.800 ;
        RECT 28.600 63.800 29.000 64.200 ;
        RECT 28.600 45.800 29.000 46.200 ;
        RECT 28.600 45.200 28.900 45.800 ;
        RECT 28.600 44.800 29.000 45.200 ;
        RECT 27.000 23.100 27.400 23.200 ;
        RECT 27.800 23.100 28.200 23.200 ;
        RECT 27.000 22.800 28.200 23.100 ;
        RECT 27.000 1.100 27.400 1.200 ;
        RECT 27.800 1.100 28.200 1.200 ;
        RECT 27.000 0.800 28.200 1.100 ;
      LAYER via3 ;
        RECT 76.600 81.800 77.000 82.200 ;
        RECT 27.800 0.800 28.200 1.200 ;
      LAYER metal4 ;
        RECT 76.600 81.800 77.000 82.200 ;
        RECT 76.600 68.200 76.900 81.800 ;
        RECT 76.600 67.800 77.000 68.200 ;
        RECT 28.600 64.800 29.000 65.200 ;
        RECT 28.600 46.200 28.900 64.800 ;
        RECT 28.600 45.800 29.000 46.200 ;
        RECT 27.000 22.800 27.400 23.200 ;
        RECT 27.000 1.100 27.300 22.800 ;
        RECT 27.800 1.100 28.200 1.200 ;
        RECT 27.000 0.800 28.200 1.100 ;
    END
  END b[3]
  PIN b[4]
    PORT
      LAYER metal1 ;
        RECT 59.000 84.400 59.400 85.200 ;
        RECT 61.400 84.400 61.800 85.200 ;
        RECT 35.800 75.800 36.200 76.600 ;
        RECT 42.600 74.800 43.400 75.200 ;
        RECT 39.800 73.800 40.200 74.600 ;
        RECT 46.200 73.800 46.600 74.600 ;
        RECT 76.600 53.400 77.000 54.200 ;
        RECT 22.200 25.800 22.600 26.200 ;
        RECT 24.200 25.800 25.000 26.200 ;
        RECT 84.600 25.800 85.000 26.600 ;
        RECT 22.200 25.200 22.500 25.800 ;
        RECT 22.200 24.400 22.600 25.200 ;
        RECT 79.800 14.800 80.200 15.600 ;
      LAYER via1 ;
        RECT 59.000 84.800 59.400 85.200 ;
        RECT 61.400 84.800 61.800 85.200 ;
        RECT 43.000 74.800 43.400 75.200 ;
        RECT 76.600 53.800 77.000 54.200 ;
        RECT 24.600 25.800 25.000 26.200 ;
      LAYER metal2 ;
        RECT 59.000 84.800 59.400 85.200 ;
        RECT 61.400 84.800 61.800 85.200 ;
        RECT 59.000 83.200 59.300 84.800 ;
        RECT 61.400 83.200 61.700 84.800 ;
        RECT 46.200 82.800 46.600 83.200 ;
        RECT 59.000 82.800 59.400 83.200 ;
        RECT 61.400 82.800 61.800 83.200 ;
        RECT 35.800 76.800 36.200 77.200 ;
        RECT 39.800 76.800 40.200 77.200 ;
        RECT 35.800 76.200 36.100 76.800 ;
        RECT 35.800 75.800 36.200 76.200 ;
        RECT 35.800 75.200 36.100 75.800 ;
        RECT 35.800 74.800 36.200 75.200 ;
        RECT 39.800 74.200 40.100 76.800 ;
        RECT 43.000 74.800 43.400 75.200 ;
        RECT 43.000 74.200 43.300 74.800 ;
        RECT 46.200 74.200 46.500 82.800 ;
        RECT 39.800 73.800 40.200 74.200 ;
        RECT 43.000 73.800 43.400 74.200 ;
        RECT 45.400 74.100 45.800 74.200 ;
        RECT 46.200 74.100 46.600 74.200 ;
        RECT 45.400 73.800 46.600 74.100 ;
        RECT 76.600 53.800 77.000 54.200 ;
        RECT 76.600 53.200 76.900 53.800 ;
        RECT 76.600 52.800 77.000 53.200 ;
        RECT 22.200 25.800 22.600 26.200 ;
        RECT 24.600 25.800 25.000 26.200 ;
        RECT 83.800 26.100 84.200 26.200 ;
        RECT 84.600 26.100 85.000 26.200 ;
        RECT 83.800 25.800 85.000 26.100 ;
        RECT 22.200 25.200 22.500 25.800 ;
        RECT 24.600 25.200 24.900 25.800 ;
        RECT 22.200 24.800 22.600 25.200 ;
        RECT 24.600 24.800 25.000 25.200 ;
        RECT 79.800 15.100 80.200 15.200 ;
        RECT 80.600 15.100 81.000 15.200 ;
        RECT 79.800 14.800 81.000 15.100 ;
        RECT 80.600 -1.800 80.900 14.800 ;
        RECT 80.600 -2.200 81.000 -1.800 ;
      LAYER via2 ;
        RECT 80.600 14.800 81.000 15.200 ;
      LAYER metal3 ;
        RECT 46.200 83.100 46.600 83.200 ;
        RECT 59.000 83.100 59.400 83.200 ;
        RECT 61.400 83.100 61.800 83.200 ;
        RECT 62.200 83.100 62.600 83.200 ;
        RECT 46.200 82.800 62.600 83.100 ;
        RECT 35.800 77.100 36.200 77.200 ;
        RECT 39.800 77.100 40.200 77.200 ;
        RECT 35.800 76.800 40.200 77.100 ;
        RECT 31.000 75.100 31.400 75.200 ;
        RECT 35.800 75.100 36.200 75.200 ;
        RECT 31.000 74.800 36.200 75.100 ;
        RECT 39.800 74.100 40.200 74.200 ;
        RECT 43.000 74.100 43.400 74.200 ;
        RECT 45.400 74.100 45.800 74.200 ;
        RECT 39.800 73.800 45.800 74.100 ;
        RECT 62.200 53.100 62.600 53.200 ;
        RECT 76.600 53.100 77.000 53.200 ;
        RECT 83.000 53.100 83.400 53.200 ;
        RECT 62.200 52.800 83.400 53.100 ;
        RECT 83.000 26.100 83.400 26.200 ;
        RECT 83.800 26.100 84.200 26.200 ;
        RECT 83.000 25.800 84.200 26.100 ;
        RECT 22.200 25.100 22.600 25.200 ;
        RECT 24.600 25.100 25.000 25.200 ;
        RECT 31.000 25.100 31.400 25.200 ;
        RECT 22.200 24.800 31.400 25.100 ;
        RECT 80.600 15.100 81.000 15.200 ;
        RECT 83.000 15.100 83.400 15.200 ;
        RECT 80.600 14.800 83.400 15.100 ;
      LAYER via3 ;
        RECT 62.200 82.800 62.600 83.200 ;
        RECT 83.000 52.800 83.400 53.200 ;
        RECT 31.000 24.800 31.400 25.200 ;
        RECT 83.000 14.800 83.400 15.200 ;
      LAYER metal4 ;
        RECT 62.200 82.800 62.600 83.200 ;
        RECT 31.000 74.800 31.400 75.200 ;
        RECT 31.000 25.200 31.300 74.800 ;
        RECT 62.200 53.200 62.500 82.800 ;
        RECT 62.200 52.800 62.600 53.200 ;
        RECT 83.000 52.800 83.400 53.200 ;
        RECT 83.000 26.200 83.300 52.800 ;
        RECT 83.000 25.800 83.400 26.200 ;
        RECT 31.000 24.800 31.400 25.200 ;
        RECT 83.000 15.200 83.300 25.800 ;
        RECT 83.000 14.800 83.400 15.200 ;
    END
  END b[4]
  PIN b[5]
    PORT
      LAYER metal1 ;
        RECT 36.600 64.400 37.000 65.200 ;
        RECT 53.400 64.400 53.800 65.200 ;
        RECT 69.400 15.100 69.800 15.200 ;
        RECT 71.000 15.100 71.400 15.200 ;
        RECT 69.400 14.800 71.400 15.100 ;
        RECT 71.000 14.400 71.400 14.800 ;
        RECT 62.200 12.400 62.600 13.200 ;
        RECT 67.000 5.400 67.400 6.200 ;
      LAYER via1 ;
        RECT 36.600 64.800 37.000 65.200 ;
        RECT 53.400 64.800 53.800 65.200 ;
        RECT 62.200 12.800 62.600 13.200 ;
        RECT 67.000 5.800 67.400 6.200 ;
      LAYER metal2 ;
        RECT 36.600 64.800 37.000 65.200 ;
        RECT 53.400 64.800 53.800 65.200 ;
        RECT 36.600 64.200 36.900 64.800 ;
        RECT 53.400 64.200 53.700 64.800 ;
        RECT 36.600 63.800 37.000 64.200 ;
        RECT 53.400 63.800 53.800 64.200 ;
        RECT 69.400 14.800 69.800 15.200 ;
        RECT 69.400 14.200 69.700 14.800 ;
        RECT 62.200 13.800 62.600 14.200 ;
        RECT 67.000 13.800 67.400 14.200 ;
        RECT 69.400 13.800 69.800 14.200 ;
        RECT 62.200 13.200 62.500 13.800 ;
        RECT 62.200 12.800 62.600 13.200 ;
        RECT 67.000 6.200 67.300 13.800 ;
        RECT 67.000 6.100 67.400 6.200 ;
        RECT 67.000 5.800 68.100 6.100 ;
        RECT 67.800 -1.800 68.100 5.800 ;
        RECT 67.800 -2.200 68.200 -1.800 ;
      LAYER metal3 ;
        RECT 36.600 64.100 37.000 64.200 ;
        RECT 53.400 64.100 53.800 64.200 ;
        RECT 59.800 64.100 60.200 64.200 ;
        RECT 36.600 63.800 60.200 64.100 ;
        RECT 59.800 14.100 60.200 14.200 ;
        RECT 62.200 14.100 62.600 14.200 ;
        RECT 67.000 14.100 67.400 14.200 ;
        RECT 69.400 14.100 69.800 14.200 ;
        RECT 59.800 13.800 69.800 14.100 ;
      LAYER via3 ;
        RECT 59.800 63.800 60.200 64.200 ;
      LAYER metal4 ;
        RECT 59.800 63.800 60.200 64.200 ;
        RECT 59.800 14.200 60.100 63.800 ;
        RECT 59.800 13.800 60.200 14.200 ;
    END
  END b[5]
  PIN b[6]
    PORT
      LAYER metal1 ;
        RECT 72.600 6.800 73.000 7.600 ;
        RECT 75.000 6.100 75.400 6.200 ;
        RECT 76.600 6.100 77.000 6.600 ;
        RECT 75.000 5.800 77.000 6.100 ;
        RECT 75.000 5.400 75.400 5.800 ;
      LAYER metal2 ;
        RECT 72.600 6.800 73.000 7.200 ;
        RECT 72.600 5.200 72.900 6.800 ;
        RECT 75.000 5.800 75.400 6.200 ;
        RECT 75.000 5.200 75.300 5.800 ;
        RECT 72.600 4.800 73.000 5.200 ;
        RECT 75.000 4.800 75.400 5.200 ;
        RECT 75.000 -1.800 75.300 4.800 ;
        RECT 75.000 -2.200 75.400 -1.800 ;
      LAYER metal3 ;
        RECT 72.600 5.100 73.000 5.200 ;
        RECT 75.000 5.100 75.400 5.200 ;
        RECT 72.600 4.800 75.400 5.100 ;
    END
  END b[6]
  PIN b[7]
    PORT
      LAYER metal1 ;
        RECT 124.600 6.100 125.000 6.200 ;
        RECT 125.400 6.100 125.800 6.200 ;
        RECT 124.600 5.800 125.800 6.100 ;
        RECT 124.600 5.400 125.000 5.800 ;
        RECT 59.000 3.800 59.400 5.200 ;
        RECT 127.000 4.400 127.400 5.200 ;
      LAYER via1 ;
        RECT 125.400 5.800 125.800 6.200 ;
        RECT 127.000 4.800 127.400 5.200 ;
      LAYER metal2 ;
        RECT 125.400 5.800 125.800 6.200 ;
        RECT 59.000 3.800 59.400 4.200 ;
        RECT 59.000 2.200 59.300 3.800 ;
        RECT 125.400 2.200 125.700 5.800 ;
        RECT 127.000 4.800 127.400 5.200 ;
        RECT 59.000 1.800 59.400 2.200 ;
        RECT 125.400 1.800 125.800 2.200 ;
        RECT 126.200 2.100 126.600 2.200 ;
        RECT 127.000 2.100 127.300 4.800 ;
        RECT 126.200 1.800 127.300 2.100 ;
        RECT 126.200 -1.800 126.500 1.800 ;
        RECT 126.200 -2.200 126.600 -1.800 ;
      LAYER metal3 ;
        RECT 59.000 2.100 59.400 2.200 ;
        RECT 125.400 2.100 125.800 2.200 ;
        RECT 126.200 2.100 126.600 2.200 ;
        RECT 59.000 1.800 126.600 2.100 ;
    END
  END b[7]
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 91.000 127.800 91.800 128.200 ;
        RECT 110.200 127.800 111.000 128.200 ;
        RECT 129.400 127.800 130.200 128.200 ;
        RECT 90.200 112.800 91.000 113.200 ;
        RECT 130.200 112.800 131.000 113.200 ;
        RECT 111.000 107.800 111.800 108.200 ;
        RECT 131.800 107.800 132.600 108.200 ;
        RECT 131.800 92.800 132.600 93.200 ;
      LAYER metal2 ;
        RECT 91.000 132.800 91.400 133.200 ;
        RECT 91.000 128.200 91.300 132.800 ;
        RECT 91.000 127.800 91.400 128.200 ;
        RECT 110.200 127.800 110.600 128.200 ;
        RECT 129.400 127.800 129.800 128.200 ;
        RECT 91.000 119.100 91.300 127.800 ;
        RECT 110.200 127.200 110.500 127.800 ;
        RECT 110.200 126.800 110.600 127.200 ;
        RECT 129.400 122.100 129.700 127.800 ;
        RECT 129.400 121.800 130.500 122.100 ;
        RECT 90.200 118.800 91.300 119.100 ;
        RECT 90.200 113.200 90.500 118.800 ;
        RECT 130.200 113.200 130.500 121.800 ;
        RECT 90.200 112.800 90.600 113.200 ;
        RECT 130.200 112.800 130.600 113.200 ;
        RECT 130.200 109.200 130.500 112.800 ;
        RECT 111.000 108.800 111.400 109.200 ;
        RECT 130.200 108.800 130.600 109.200 ;
        RECT 131.800 108.800 132.200 109.200 ;
        RECT 111.000 108.200 111.300 108.800 ;
        RECT 131.800 108.200 132.100 108.800 ;
        RECT 111.000 107.800 111.400 108.200 ;
        RECT 131.800 107.800 132.200 108.200 ;
        RECT 131.800 93.200 132.100 107.800 ;
        RECT 131.800 92.800 132.200 93.200 ;
      LAYER metal3 ;
        RECT 91.000 128.100 91.400 128.200 ;
        RECT 110.200 128.100 110.600 128.200 ;
        RECT 91.000 127.800 110.600 128.100 ;
        RECT 110.200 127.200 110.500 127.800 ;
        RECT 110.200 126.800 110.600 127.200 ;
        RECT 110.200 109.100 110.600 109.200 ;
        RECT 111.000 109.100 111.400 109.200 ;
        RECT 130.200 109.100 130.600 109.200 ;
        RECT 131.800 109.100 132.200 109.200 ;
        RECT 110.200 108.800 132.200 109.100 ;
      LAYER via3 ;
        RECT 110.200 127.800 110.600 128.200 ;
      LAYER metal4 ;
        RECT 110.200 127.800 110.600 128.200 ;
        RECT 110.200 109.200 110.500 127.800 ;
        RECT 110.200 108.800 110.600 109.200 ;
    END
  END clk
  PIN rst
    PORT
      LAYER metal1 ;
        RECT 79.000 126.800 79.400 127.600 ;
      LAYER metal2 ;
        RECT 77.400 132.800 77.800 133.200 ;
        RECT 77.400 128.200 77.700 132.800 ;
        RECT 77.400 127.800 77.800 128.200 ;
        RECT 79.000 127.800 79.400 128.200 ;
        RECT 79.000 127.200 79.300 127.800 ;
        RECT 79.000 126.800 79.400 127.200 ;
      LAYER metal3 ;
        RECT 77.400 128.100 77.800 128.200 ;
        RECT 79.000 128.100 79.400 128.200 ;
        RECT 77.400 127.800 79.400 128.100 ;
    END
  END rst
  PIN en
    PORT
      LAYER metal1 ;
        RECT 103.800 113.400 104.200 114.200 ;
        RECT 94.200 105.400 94.600 106.200 ;
        RECT 96.600 105.400 97.000 106.200 ;
        RECT 122.200 106.100 122.600 106.600 ;
        RECT 123.000 106.100 123.400 106.200 ;
        RECT 122.200 105.800 123.400 106.100 ;
        RECT 117.000 96.800 117.400 97.200 ;
        RECT 117.100 96.200 117.400 96.800 ;
        RECT 117.100 95.900 117.800 96.200 ;
        RECT 117.400 95.800 117.800 95.900 ;
        RECT 123.000 94.800 123.400 95.600 ;
        RECT 143.000 85.800 143.400 86.600 ;
        RECT 140.200 76.800 140.600 77.200 ;
        RECT 140.200 76.200 140.500 76.800 ;
        RECT 139.800 75.900 140.500 76.200 ;
        RECT 139.800 75.800 140.200 75.900 ;
        RECT 129.000 56.800 129.400 57.200 ;
        RECT 129.100 56.200 129.400 56.800 ;
        RECT 129.100 55.900 129.800 56.200 ;
        RECT 129.400 55.800 129.800 55.900 ;
        RECT 127.000 45.100 127.400 45.200 ;
        RECT 127.000 44.800 127.700 45.100 ;
        RECT 127.400 44.200 127.700 44.800 ;
        RECT 127.400 43.800 127.800 44.200 ;
        RECT 130.600 16.800 131.000 17.200 ;
        RECT 130.700 16.200 131.000 16.800 ;
        RECT 130.700 15.900 131.400 16.200 ;
        RECT 131.000 15.800 131.400 15.900 ;
        RECT 88.600 5.800 89.000 6.200 ;
        RECT 88.600 5.200 88.900 5.800 ;
        RECT 88.600 5.100 89.000 5.200 ;
        RECT 103.000 5.100 103.400 5.200 ;
        RECT 88.600 4.800 89.300 5.100 ;
        RECT 89.000 4.200 89.300 4.800 ;
        RECT 102.700 4.800 103.400 5.100 ;
        RECT 119.800 5.100 120.200 5.200 ;
        RECT 119.800 4.800 120.500 5.100 ;
        RECT 102.700 4.200 103.000 4.800 ;
        RECT 89.000 3.800 89.400 4.200 ;
        RECT 102.600 3.800 103.000 4.200 ;
        RECT 120.200 4.200 120.500 4.800 ;
        RECT 120.200 3.800 120.600 4.200 ;
      LAYER via1 ;
        RECT 103.800 113.800 104.200 114.200 ;
        RECT 94.200 105.800 94.600 106.200 ;
        RECT 96.600 105.800 97.000 106.200 ;
        RECT 123.000 105.800 123.400 106.200 ;
        RECT 103.000 4.800 103.400 5.200 ;
      LAYER metal2 ;
        RECT 103.800 113.800 104.200 114.200 ;
        RECT 103.800 106.200 104.100 113.800 ;
        RECT 94.200 106.100 94.600 106.200 ;
        RECT 95.000 106.100 95.400 106.200 ;
        RECT 94.200 105.800 95.400 106.100 ;
        RECT 96.600 106.100 97.000 106.200 ;
        RECT 97.400 106.100 97.800 106.200 ;
        RECT 96.600 105.800 97.800 106.100 ;
        RECT 103.800 105.800 104.200 106.200 ;
        RECT 123.000 105.800 123.400 106.200 ;
        RECT 117.400 95.800 117.800 96.200 ;
        RECT 117.400 91.200 117.700 95.800 ;
        RECT 123.000 95.200 123.300 105.800 ;
        RECT 123.000 94.800 123.400 95.200 ;
        RECT 123.000 91.200 123.300 94.800 ;
        RECT 117.400 90.800 117.800 91.200 ;
        RECT 123.000 90.800 123.400 91.200 ;
        RECT 142.200 90.800 142.600 91.200 ;
        RECT 142.200 86.200 142.500 90.800 ;
        RECT 139.800 85.800 140.200 86.200 ;
        RECT 142.200 86.100 142.600 86.200 ;
        RECT 143.000 86.100 143.400 86.200 ;
        RECT 142.200 85.800 143.400 86.100 ;
        RECT 139.800 76.200 140.100 85.800 ;
        RECT 139.800 75.800 140.200 76.200 ;
        RECT 139.800 70.200 140.100 75.800 ;
        RECT 129.400 69.800 129.800 70.200 ;
        RECT 139.800 69.800 140.200 70.200 ;
        RECT 129.400 56.200 129.700 69.800 ;
        RECT 129.400 55.800 129.800 56.200 ;
        RECT 129.400 55.200 129.700 55.800 ;
        RECT 129.400 54.800 129.800 55.200 ;
        RECT 127.000 44.800 127.400 45.200 ;
        RECT 127.000 44.200 127.300 44.800 ;
        RECT 127.000 43.800 127.400 44.200 ;
        RECT 130.200 16.100 130.600 16.200 ;
        RECT 131.000 16.100 131.400 16.200 ;
        RECT 130.200 15.800 131.400 16.100 ;
        RECT 88.600 5.800 89.000 6.200 ;
        RECT 88.600 5.200 88.900 5.800 ;
        RECT 88.600 4.800 89.000 5.200 ;
        RECT 102.200 5.100 102.600 5.200 ;
        RECT 103.000 5.100 103.400 5.200 ;
        RECT 102.200 4.800 103.400 5.100 ;
        RECT 119.000 5.100 119.400 5.200 ;
        RECT 119.800 5.100 120.200 5.200 ;
        RECT 119.000 4.800 120.200 5.100 ;
        RECT 120.600 4.800 121.000 5.200 ;
        RECT 120.600 -1.800 120.900 4.800 ;
        RECT 120.600 -2.200 121.000 -1.800 ;
      LAYER via2 ;
        RECT 95.000 105.800 95.400 106.200 ;
        RECT 97.400 105.800 97.800 106.200 ;
      LAYER metal3 ;
        RECT 95.000 106.100 95.400 106.200 ;
        RECT 97.400 106.100 97.800 106.200 ;
        RECT 103.800 106.100 104.200 106.200 ;
        RECT 123.000 106.100 123.400 106.200 ;
        RECT 95.000 105.800 123.400 106.100 ;
        RECT 117.400 91.100 117.800 91.200 ;
        RECT 123.000 91.100 123.400 91.200 ;
        RECT 142.200 91.100 142.600 91.200 ;
        RECT 117.400 90.800 142.600 91.100 ;
        RECT 139.800 86.100 140.200 86.200 ;
        RECT 142.200 86.100 142.600 86.200 ;
        RECT 139.800 85.800 142.600 86.100 ;
        RECT 129.400 70.100 129.800 70.200 ;
        RECT 139.800 70.100 140.200 70.200 ;
        RECT 129.400 69.800 140.200 70.100 ;
        RECT 129.400 55.800 129.800 56.200 ;
        RECT 129.400 55.200 129.700 55.800 ;
        RECT 129.400 54.800 129.800 55.200 ;
        RECT 127.000 44.100 127.400 44.200 ;
        RECT 129.400 44.100 129.800 44.200 ;
        RECT 127.000 43.800 129.800 44.100 ;
        RECT 129.400 16.100 129.800 16.200 ;
        RECT 130.200 16.100 130.600 16.200 ;
        RECT 129.400 15.800 130.600 16.100 ;
        RECT 88.600 5.100 89.000 5.200 ;
        RECT 102.200 5.100 102.600 5.200 ;
        RECT 119.000 5.100 119.400 5.200 ;
        RECT 120.600 5.100 121.000 5.200 ;
        RECT 130.200 5.100 130.600 5.200 ;
        RECT 88.600 4.800 130.600 5.100 ;
      LAYER via3 ;
        RECT 129.400 43.800 129.800 44.200 ;
        RECT 130.200 4.800 130.600 5.200 ;
      LAYER metal4 ;
        RECT 129.400 55.800 129.800 56.200 ;
        RECT 129.400 44.200 129.700 55.800 ;
        RECT 129.400 43.800 129.800 44.200 ;
        RECT 129.400 16.200 129.700 43.800 ;
        RECT 129.400 16.100 129.800 16.200 ;
        RECT 129.400 15.800 130.500 16.100 ;
        RECT 130.200 5.200 130.500 15.800 ;
        RECT 130.200 4.800 130.600 5.200 ;
    END
  END en
  PIN opcode[0]
    PORT
      LAYER metal1 ;
        RECT 149.400 126.800 149.800 127.600 ;
        RECT 148.600 47.800 149.000 48.600 ;
        RECT 143.800 35.800 144.200 36.600 ;
        RECT 147.600 34.200 148.000 34.600 ;
        RECT 147.700 34.100 148.200 34.200 ;
        RECT 148.600 34.100 149.000 34.200 ;
        RECT 147.700 33.800 149.000 34.100 ;
      LAYER via1 ;
        RECT 148.600 33.800 149.000 34.200 ;
      LAYER metal2 ;
        RECT 151.800 132.100 152.200 132.200 ;
        RECT 150.200 131.800 152.200 132.100 ;
        RECT 149.400 127.100 149.800 127.200 ;
        RECT 150.200 127.100 150.500 131.800 ;
        RECT 149.400 126.800 150.500 127.100 ;
        RECT 149.400 120.200 149.700 126.800 ;
        RECT 149.400 119.800 149.800 120.200 ;
        RECT 148.600 51.800 149.000 52.200 ;
        RECT 148.600 48.200 148.900 51.800 ;
        RECT 148.600 47.800 149.000 48.200 ;
        RECT 148.600 37.200 148.900 47.800 ;
        RECT 143.800 36.800 144.200 37.200 ;
        RECT 148.600 36.800 149.000 37.200 ;
        RECT 143.800 36.200 144.100 36.800 ;
        RECT 143.800 35.800 144.200 36.200 ;
        RECT 148.600 34.200 148.900 36.800 ;
        RECT 148.600 33.800 149.000 34.200 ;
      LAYER via2 ;
        RECT 151.800 131.800 152.200 132.200 ;
      LAYER metal3 ;
        RECT 151.800 132.100 152.200 132.200 ;
        RECT 153.400 132.100 153.800 132.200 ;
        RECT 151.800 131.800 153.800 132.100 ;
        RECT 149.400 119.800 149.800 120.200 ;
        RECT 149.400 119.200 149.700 119.800 ;
        RECT 149.400 118.800 149.800 119.200 ;
        RECT 148.600 52.100 149.000 52.200 ;
        RECT 149.400 52.100 149.800 52.200 ;
        RECT 148.600 51.800 149.800 52.100 ;
        RECT 143.800 37.100 144.200 37.200 ;
        RECT 148.600 37.100 149.000 37.200 ;
        RECT 143.800 36.800 149.000 37.100 ;
      LAYER via3 ;
        RECT 149.400 51.800 149.800 52.200 ;
      LAYER metal4 ;
        RECT 149.400 118.800 149.800 119.200 ;
        RECT 149.400 52.200 149.700 118.800 ;
        RECT 149.400 51.800 149.800 52.200 ;
    END
  END opcode[0]
  PIN opcode[1]
    PORT
      LAYER metal1 ;
        RECT 145.400 33.400 145.800 34.200 ;
        RECT 148.600 32.400 149.000 33.200 ;
        RECT 148.600 27.800 149.000 28.600 ;
      LAYER via1 ;
        RECT 145.400 33.800 145.800 34.200 ;
        RECT 148.600 32.800 149.000 33.200 ;
      LAYER metal2 ;
        RECT 145.400 33.800 145.800 34.200 ;
        RECT 145.400 32.200 145.700 33.800 ;
        RECT 148.600 32.800 149.000 33.200 ;
        RECT 148.600 32.200 148.900 32.800 ;
        RECT 145.400 31.800 145.800 32.200 ;
        RECT 148.600 31.800 149.000 32.200 ;
        RECT 148.600 28.200 148.900 31.800 ;
        RECT 148.600 27.800 149.000 28.200 ;
      LAYER metal3 ;
        RECT 145.400 32.100 145.800 32.200 ;
        RECT 148.600 32.100 149.000 32.200 ;
        RECT 145.400 31.800 149.000 32.100 ;
        RECT 148.600 28.100 149.000 28.200 ;
        RECT 153.400 28.100 153.800 28.200 ;
        RECT 148.600 27.800 153.800 28.100 ;
    END
  END opcode[1]
  PIN opcode[2]
    PORT
      LAYER metal1 ;
        RECT 146.200 126.800 146.600 127.600 ;
        RECT 146.200 52.400 146.600 53.200 ;
        RECT 143.000 32.400 143.400 33.200 ;
        RECT 143.800 27.800 144.200 28.600 ;
        RECT 149.400 13.100 149.800 13.200 ;
        RECT 150.200 13.100 150.600 13.200 ;
        RECT 149.400 12.800 150.600 13.100 ;
        RECT 149.400 12.400 149.800 12.800 ;
      LAYER via1 ;
        RECT 146.200 52.800 146.600 53.200 ;
        RECT 143.000 32.800 143.400 33.200 ;
        RECT 150.200 12.800 150.600 13.200 ;
      LAYER metal2 ;
        RECT 146.200 126.800 146.600 127.200 ;
        RECT 146.200 117.200 146.500 126.800 ;
        RECT 146.200 116.800 146.600 117.200 ;
        RECT 146.200 53.800 146.600 54.200 ;
        RECT 146.200 53.200 146.500 53.800 ;
        RECT 146.200 52.800 146.600 53.200 ;
        RECT 143.000 33.100 143.400 33.200 ;
        RECT 143.800 33.100 144.200 33.200 ;
        RECT 143.000 32.800 144.200 33.100 ;
        RECT 143.800 28.200 144.100 32.800 ;
        RECT 143.800 27.800 144.200 28.200 ;
        RECT 143.800 26.200 144.100 27.800 ;
        RECT 143.800 25.800 144.200 26.200 ;
        RECT 150.200 25.800 150.600 26.200 ;
        RECT 150.200 13.200 150.500 25.800 ;
        RECT 150.200 12.800 150.600 13.200 ;
      LAYER via2 ;
        RECT 143.800 32.800 144.200 33.200 ;
      LAYER metal3 ;
        RECT 146.200 116.800 146.600 117.200 ;
        RECT 146.200 116.200 146.500 116.800 ;
        RECT 146.200 115.800 146.600 116.200 ;
        RECT 146.200 53.800 146.600 54.200 ;
        RECT 146.200 53.200 146.500 53.800 ;
        RECT 146.200 52.800 146.600 53.200 ;
        RECT 143.800 33.100 144.200 33.200 ;
        RECT 146.200 33.100 146.600 33.200 ;
        RECT 143.800 32.800 146.600 33.100 ;
        RECT 143.800 26.100 144.200 26.200 ;
        RECT 150.200 26.100 150.600 26.200 ;
        RECT 153.400 26.100 153.800 26.200 ;
        RECT 143.800 25.800 153.800 26.100 ;
      LAYER via3 ;
        RECT 146.200 32.800 146.600 33.200 ;
      LAYER metal4 ;
        RECT 146.200 115.800 146.600 116.200 ;
        RECT 146.200 53.200 146.500 115.800 ;
        RECT 146.200 52.800 146.600 53.200 ;
        RECT 146.200 33.200 146.500 52.800 ;
        RECT 146.200 32.800 146.600 33.200 ;
    END
  END opcode[2]
  PIN out[0]
    PORT
      LAYER metal1 ;
        RECT 147.800 86.200 148.200 89.900 ;
        RECT 147.900 85.100 148.200 86.200 ;
        RECT 147.800 81.100 148.200 85.100 ;
      LAYER via1 ;
        RECT 147.800 83.800 148.200 84.200 ;
      LAYER metal2 ;
        RECT 147.800 84.800 148.200 85.200 ;
        RECT 147.800 84.200 148.100 84.800 ;
        RECT 147.800 83.800 148.200 84.200 ;
      LAYER metal3 ;
        RECT 147.800 85.100 148.200 85.200 ;
        RECT 153.400 85.100 153.800 85.200 ;
        RECT 147.800 84.800 153.800 85.100 ;
    END
  END out[0]
  PIN out[1]
    PORT
      LAYER metal1 ;
        RECT 147.800 95.900 148.200 99.900 ;
        RECT 147.900 94.800 148.200 95.900 ;
        RECT 147.800 91.100 148.200 94.800 ;
      LAYER via1 ;
        RECT 147.800 96.800 148.200 97.200 ;
      LAYER metal2 ;
        RECT 147.800 96.800 148.200 97.200 ;
        RECT 147.800 96.200 148.100 96.800 ;
        RECT 147.800 95.800 148.200 96.200 ;
      LAYER metal3 ;
        RECT 147.800 96.100 148.200 96.200 ;
        RECT 147.800 95.800 151.300 96.100 ;
        RECT 151.000 95.100 151.300 95.800 ;
        RECT 153.400 95.100 153.800 95.200 ;
        RECT 151.000 94.800 153.800 95.100 ;
    END
  END out[1]
  PIN out[2]
    PORT
      LAYER metal1 ;
        RECT 143.000 95.900 143.400 99.900 ;
        RECT 143.100 94.800 143.400 95.900 ;
        RECT 143.000 91.100 143.400 94.800 ;
      LAYER via1 ;
        RECT 143.000 96.800 143.400 97.200 ;
      LAYER metal2 ;
        RECT 143.000 97.100 143.400 97.200 ;
        RECT 143.800 97.100 144.200 97.200 ;
        RECT 143.000 96.800 144.200 97.100 ;
      LAYER via2 ;
        RECT 143.800 96.800 144.200 97.200 ;
      LAYER metal3 ;
        RECT 143.800 97.100 144.200 97.200 ;
        RECT 153.400 97.100 153.800 97.200 ;
        RECT 143.000 96.800 153.800 97.100 ;
    END
  END out[2]
  PIN out[3]
    PORT
      LAYER metal1 ;
        RECT 145.400 115.900 145.800 119.900 ;
        RECT 145.500 114.800 145.800 115.900 ;
        RECT 145.400 111.100 145.800 114.800 ;
      LAYER via1 ;
        RECT 145.400 113.800 145.800 114.200 ;
      LAYER metal2 ;
        RECT 145.400 114.800 145.800 115.200 ;
        RECT 145.400 114.200 145.700 114.800 ;
        RECT 145.400 113.800 145.800 114.200 ;
      LAYER metal3 ;
        RECT 145.400 115.100 145.800 115.200 ;
        RECT 153.400 115.100 153.800 115.200 ;
        RECT 145.400 114.800 153.800 115.100 ;
    END
  END out[3]
  PIN out[4]
    PORT
      LAYER metal1 ;
        RECT 143.000 115.900 143.400 119.900 ;
        RECT 143.100 114.800 143.400 115.900 ;
        RECT 143.000 111.100 143.400 114.800 ;
      LAYER via1 ;
        RECT 143.000 117.800 143.400 118.200 ;
      LAYER metal2 ;
        RECT 143.000 118.800 143.400 119.200 ;
        RECT 143.000 118.200 143.300 118.800 ;
        RECT 143.000 117.800 143.400 118.200 ;
      LAYER metal3 ;
        RECT 143.000 118.800 143.400 119.200 ;
        RECT 143.000 118.100 143.300 118.800 ;
        RECT 143.000 117.800 153.700 118.100 ;
        RECT 153.400 117.200 153.700 117.800 ;
        RECT 153.400 116.800 153.800 117.200 ;
    END
  END out[4]
  PIN out[5]
    PORT
      LAYER metal1 ;
        RECT 140.600 126.200 141.000 129.900 ;
        RECT 140.700 125.100 141.000 126.200 ;
        RECT 140.600 121.100 141.000 125.100 ;
      LAYER via1 ;
        RECT 140.600 122.800 141.000 123.200 ;
      LAYER metal2 ;
        RECT 140.600 123.800 141.000 124.200 ;
        RECT 140.600 123.200 140.900 123.800 ;
        RECT 140.600 122.800 141.000 123.200 ;
      LAYER metal3 ;
        RECT 140.600 123.800 141.000 124.200 ;
        RECT 153.400 123.800 153.800 124.200 ;
        RECT 140.600 123.100 140.900 123.800 ;
        RECT 153.400 123.100 153.700 123.800 ;
        RECT 140.600 122.800 153.700 123.100 ;
    END
  END out[5]
  PIN out[6]
    PORT
      LAYER metal1 ;
        RECT 143.000 126.200 143.400 129.900 ;
        RECT 143.100 125.100 143.400 126.200 ;
        RECT 143.000 121.100 143.400 125.100 ;
      LAYER via1 ;
        RECT 143.000 126.800 143.400 127.200 ;
      LAYER metal2 ;
        RECT 143.000 126.800 143.400 127.200 ;
        RECT 143.000 126.200 143.300 126.800 ;
        RECT 143.000 125.800 143.400 126.200 ;
      LAYER metal3 ;
        RECT 143.000 126.100 143.400 126.200 ;
        RECT 153.400 126.100 153.800 126.200 ;
        RECT 143.000 125.800 153.800 126.100 ;
    END
  END out[6]
  PIN out[7]
    PORT
      LAYER metal1 ;
        RECT 145.400 126.200 145.800 129.900 ;
        RECT 145.500 125.100 145.800 126.200 ;
        RECT 145.400 121.100 145.800 125.100 ;
      LAYER via1 ;
        RECT 145.400 127.800 145.800 128.200 ;
      LAYER metal2 ;
        RECT 145.400 127.800 145.800 128.200 ;
        RECT 145.400 127.200 145.700 127.800 ;
        RECT 145.400 126.800 145.800 127.200 ;
      LAYER metal3 ;
        RECT 153.400 128.100 153.800 128.200 ;
        RECT 145.400 127.800 153.800 128.100 ;
        RECT 145.400 127.200 145.700 127.800 ;
        RECT 145.400 126.800 145.800 127.200 ;
    END
  END out[7]
  PIN zero
    PORT
      LAYER metal1 ;
        RECT 147.800 115.900 148.200 119.900 ;
        RECT 147.900 114.800 148.200 115.900 ;
        RECT 147.800 111.100 148.200 114.800 ;
      LAYER via1 ;
        RECT 147.800 118.800 148.200 119.200 ;
      LAYER metal2 ;
        RECT 148.600 129.800 149.000 130.200 ;
        RECT 148.600 123.100 148.900 129.800 ;
        RECT 147.800 122.800 148.900 123.100 ;
        RECT 147.800 119.200 148.100 122.800 ;
        RECT 147.800 118.800 148.200 119.200 ;
      LAYER metal3 ;
        RECT 148.600 130.100 149.000 130.200 ;
        RECT 153.400 130.100 153.800 130.200 ;
        RECT 148.600 129.800 153.800 130.100 ;
    END
  END zero
  OBS
      LAYER metal1 ;
        RECT 1.200 127.100 1.600 129.900 ;
        RECT 5.400 127.900 5.800 129.900 ;
        RECT 6.100 128.200 6.500 128.600 ;
        RECT 7.100 128.200 7.500 128.600 ;
        RECT 0.700 126.900 1.600 127.100 ;
        RECT 0.700 126.800 1.500 126.900 ;
        RECT 0.700 126.200 1.000 126.800 ;
        RECT 4.600 126.400 5.000 127.200 ;
        RECT 5.400 127.100 5.700 127.900 ;
        RECT 6.200 127.800 6.600 128.200 ;
        RECT 7.000 127.800 7.400 128.200 ;
        RECT 7.800 127.900 8.200 129.900 ;
        RECT 7.000 127.200 7.300 127.800 ;
        RECT 7.000 127.100 7.400 127.200 ;
        RECT 5.400 126.800 7.400 127.100 ;
        RECT 0.600 125.800 1.000 126.200 ;
        RECT 1.800 125.800 2.600 126.200 ;
        RECT 3.800 126.100 4.200 126.200 ;
        RECT 5.400 126.100 5.700 126.800 ;
        RECT 6.200 126.100 6.600 126.200 ;
        RECT 3.800 125.800 4.600 126.100 ;
        RECT 5.400 125.800 6.600 126.100 ;
        RECT 7.000 126.100 7.400 126.200 ;
        RECT 7.900 126.100 8.200 127.900 ;
        RECT 8.600 126.400 9.000 127.200 ;
        RECT 9.400 126.800 9.800 127.200 ;
        RECT 12.000 127.100 12.400 129.900 ;
        RECT 13.400 128.000 13.800 129.900 ;
        RECT 15.000 128.000 15.400 129.900 ;
        RECT 13.400 127.900 15.400 128.000 ;
        RECT 15.800 127.900 16.200 129.900 ;
        RECT 13.500 127.700 15.300 127.900 ;
        RECT 13.800 127.200 14.200 127.400 ;
        RECT 15.800 127.200 16.100 127.900 ;
        RECT 12.000 126.900 12.900 127.100 ;
        RECT 12.100 126.800 12.900 126.900 ;
        RECT 13.400 126.900 14.200 127.200 ;
        RECT 13.400 126.800 13.800 126.900 ;
        RECT 14.900 126.800 16.200 127.200 ;
        RECT 17.200 127.100 17.600 129.900 ;
        RECT 19.800 128.000 20.200 129.900 ;
        RECT 21.400 128.000 21.800 129.900 ;
        RECT 19.800 127.900 21.800 128.000 ;
        RECT 22.200 127.900 22.600 129.900 ;
        RECT 19.900 127.700 21.700 127.900 ;
        RECT 20.200 127.200 20.600 127.400 ;
        RECT 22.200 127.200 22.500 127.900 ;
        RECT 16.700 126.900 17.600 127.100 ;
        RECT 19.800 126.900 20.600 127.200 ;
        RECT 16.700 126.800 17.500 126.900 ;
        RECT 19.800 126.800 20.200 126.900 ;
        RECT 21.300 126.800 22.600 127.200 ;
        RECT 24.800 127.100 25.200 129.900 ;
        RECT 27.500 127.900 28.300 129.900 ;
        RECT 31.000 128.900 31.400 129.900 ;
        RECT 34.200 129.200 34.600 129.900 ;
        RECT 34.200 128.900 34.700 129.200 ;
        RECT 27.800 127.200 28.100 127.900 ;
        RECT 31.000 127.200 31.300 128.900 ;
        RECT 34.400 128.800 34.700 128.900 ;
        RECT 35.800 128.900 36.200 129.900 ;
        RECT 35.800 128.800 36.400 128.900 ;
        RECT 31.800 128.100 32.200 128.600 ;
        RECT 34.400 128.500 36.400 128.800 ;
        RECT 33.400 128.100 34.300 128.200 ;
        RECT 31.800 127.800 34.300 128.100 ;
        RECT 24.800 126.900 25.700 127.100 ;
        RECT 24.900 126.800 25.700 126.900 ;
        RECT 27.000 126.800 27.400 127.200 ;
        RECT 9.400 126.200 9.700 126.800 ;
        RECT 9.400 126.100 9.800 126.200 ;
        RECT 7.000 125.800 8.200 126.100 ;
        RECT 9.000 125.800 9.800 126.100 ;
        RECT 11.000 125.800 11.800 126.200 ;
        RECT 0.700 125.200 1.000 125.800 ;
        RECT 4.200 125.600 4.600 125.800 ;
        RECT 0.600 124.800 1.000 125.200 ;
        RECT 3.000 124.800 3.400 125.600 ;
        RECT 6.200 125.100 6.500 125.800 ;
        RECT 7.100 125.100 7.400 125.800 ;
        RECT 9.000 125.600 9.400 125.800 ;
        RECT 3.800 124.800 5.800 125.100 ;
        RECT 0.700 123.500 1.000 124.800 ;
        RECT 1.400 123.800 1.800 124.600 ;
        RECT 0.700 123.200 2.500 123.500 ;
        RECT 0.700 123.100 1.000 123.200 ;
        RECT 0.600 121.100 1.000 123.100 ;
        RECT 2.200 123.100 2.500 123.200 ;
        RECT 2.200 121.100 2.600 123.100 ;
        RECT 3.800 121.100 4.200 124.800 ;
        RECT 5.400 121.100 5.800 124.800 ;
        RECT 6.200 121.100 6.600 125.100 ;
        RECT 7.000 121.100 7.400 125.100 ;
        RECT 7.800 124.800 9.800 125.100 ;
        RECT 10.200 124.800 10.600 125.600 ;
        RECT 12.600 125.200 12.900 126.800 ;
        RECT 14.200 125.800 14.600 126.600 ;
        RECT 12.600 124.800 13.000 125.200 ;
        RECT 14.900 125.100 15.200 126.800 ;
        RECT 16.700 125.200 17.000 126.800 ;
        RECT 17.800 125.800 18.600 126.200 ;
        RECT 19.800 126.100 20.200 126.200 ;
        RECT 20.600 126.100 21.000 126.600 ;
        RECT 19.800 125.800 21.000 126.100 ;
        RECT 15.800 125.100 16.200 125.200 ;
        RECT 14.700 124.800 15.200 125.100 ;
        RECT 15.500 124.800 16.200 125.100 ;
        RECT 16.600 124.800 17.000 125.200 ;
        RECT 19.000 124.800 19.400 125.600 ;
        RECT 21.300 125.100 21.600 126.800 ;
        RECT 23.800 125.800 24.600 126.200 ;
        RECT 22.200 125.100 22.600 125.200 ;
        RECT 21.100 124.800 21.600 125.100 ;
        RECT 21.900 124.800 22.600 125.100 ;
        RECT 23.000 125.100 23.400 125.600 ;
        RECT 25.400 125.200 25.700 126.800 ;
        RECT 27.100 126.600 27.400 126.800 ;
        RECT 27.800 126.800 28.200 127.200 ;
        RECT 28.600 127.100 29.000 127.200 ;
        RECT 31.000 127.100 31.400 127.200 ;
        RECT 28.600 126.800 31.400 127.100 ;
        RECT 34.200 126.800 35.000 127.200 ;
        RECT 27.100 126.200 27.500 126.600 ;
        RECT 27.800 126.200 28.100 126.800 ;
        RECT 28.600 126.400 29.000 126.800 ;
        RECT 26.200 125.400 26.600 126.200 ;
        RECT 27.800 125.800 28.200 126.200 ;
        RECT 29.400 126.100 29.800 126.200 ;
        RECT 29.000 125.800 29.800 126.100 ;
        RECT 27.800 125.700 28.100 125.800 ;
        RECT 27.100 125.400 28.100 125.700 ;
        RECT 29.000 125.600 29.400 125.800 ;
        RECT 30.200 125.400 30.600 126.200 ;
        RECT 23.800 125.100 24.200 125.200 ;
        RECT 23.000 124.800 24.200 125.100 ;
        RECT 25.400 124.800 25.800 125.200 ;
        RECT 27.100 125.100 27.400 125.400 ;
        RECT 31.000 125.100 31.300 126.800 ;
        RECT 35.000 125.800 35.800 126.200 ;
        RECT 36.100 125.300 36.400 128.500 ;
        RECT 39.600 127.100 40.000 129.900 ;
        RECT 42.200 128.000 42.600 129.900 ;
        RECT 43.800 128.000 44.200 129.900 ;
        RECT 42.200 127.900 44.200 128.000 ;
        RECT 44.600 127.900 45.000 129.900 ;
        RECT 47.000 127.900 47.400 129.900 ;
        RECT 47.700 128.200 48.100 128.600 ;
        RECT 42.300 127.700 44.100 127.900 ;
        RECT 42.600 127.200 43.000 127.400 ;
        RECT 44.600 127.200 44.900 127.900 ;
        RECT 39.100 126.900 40.000 127.100 ;
        RECT 42.200 126.900 43.000 127.200 ;
        RECT 43.700 127.100 45.000 127.200 ;
        RECT 46.200 127.100 46.600 127.200 ;
        RECT 39.100 126.800 39.900 126.900 ;
        RECT 42.200 126.800 42.600 126.900 ;
        RECT 43.700 126.800 46.600 127.100 ;
        RECT 36.100 125.200 37.000 125.300 ;
        RECT 39.100 125.200 39.400 126.800 ;
        RECT 40.200 125.800 41.000 126.200 ;
        RECT 43.000 125.800 43.400 126.600 ;
        RECT 7.800 121.100 8.200 124.800 ;
        RECT 9.400 121.100 9.800 124.800 ;
        RECT 11.800 123.800 12.200 124.600 ;
        RECT 12.600 123.500 12.900 124.800 ;
        RECT 11.100 123.200 12.900 123.500 ;
        RECT 11.100 123.100 11.400 123.200 ;
        RECT 11.000 121.100 11.400 123.100 ;
        RECT 12.600 123.100 12.900 123.200 ;
        RECT 12.600 121.100 13.000 123.100 ;
        RECT 14.700 121.100 15.100 124.800 ;
        RECT 15.500 124.200 15.800 124.800 ;
        RECT 15.400 123.800 15.800 124.200 ;
        RECT 16.700 123.500 17.000 124.800 ;
        RECT 17.400 123.800 17.800 124.600 ;
        RECT 16.700 123.200 18.500 123.500 ;
        RECT 16.700 123.100 17.000 123.200 ;
        RECT 16.600 121.100 17.000 123.100 ;
        RECT 18.200 123.100 18.500 123.200 ;
        RECT 18.200 121.100 18.600 123.100 ;
        RECT 21.100 122.200 21.500 124.800 ;
        RECT 21.900 124.200 22.200 124.800 ;
        RECT 21.800 124.100 22.600 124.200 ;
        RECT 21.800 123.800 24.100 124.100 ;
        RECT 24.600 123.800 25.000 124.600 ;
        RECT 20.600 121.800 21.500 122.200 ;
        RECT 21.100 121.100 21.500 121.800 ;
        RECT 23.800 123.500 24.100 123.800 ;
        RECT 25.400 123.500 25.700 124.800 ;
        RECT 23.800 123.200 25.700 123.500 ;
        RECT 23.800 121.100 24.200 123.200 ;
        RECT 25.400 123.100 25.700 123.200 ;
        RECT 25.400 121.100 25.800 123.100 ;
        RECT 26.200 121.400 26.600 125.100 ;
        RECT 27.000 121.700 27.400 125.100 ;
        RECT 27.800 124.800 29.800 125.100 ;
        RECT 27.800 121.400 28.200 124.800 ;
        RECT 26.200 121.100 28.200 121.400 ;
        RECT 29.400 121.100 29.800 124.800 ;
        RECT 30.500 124.700 31.400 125.100 ;
        RECT 36.100 124.900 37.800 125.200 ;
        RECT 37.400 124.800 37.800 124.900 ;
        RECT 39.000 124.800 39.400 125.200 ;
        RECT 41.400 124.800 41.800 125.600 ;
        RECT 43.700 125.100 44.000 126.800 ;
        RECT 46.200 126.400 46.600 126.800 ;
        RECT 45.400 126.100 45.800 126.200 ;
        RECT 47.000 126.100 47.300 127.900 ;
        RECT 47.800 127.800 48.200 128.200 ;
        RECT 52.000 127.100 52.400 129.900 ;
        RECT 54.000 127.100 54.400 129.900 ;
        RECT 59.000 128.900 59.400 129.900 ;
        RECT 60.600 129.200 61.000 129.900 ;
        RECT 58.800 128.800 59.400 128.900 ;
        RECT 60.500 128.900 61.000 129.200 ;
        RECT 60.500 128.800 60.800 128.900 ;
        RECT 58.800 128.500 60.800 128.800 ;
        RECT 57.400 128.100 57.800 128.200 ;
        RECT 58.800 128.100 59.100 128.500 ;
        RECT 57.400 127.800 59.100 128.100 ;
        RECT 60.900 127.800 61.800 128.200 ;
        RECT 63.000 128.000 63.400 129.900 ;
        RECT 64.600 128.000 65.000 129.900 ;
        RECT 63.000 127.900 65.000 128.000 ;
        RECT 65.400 127.900 65.800 129.900 ;
        RECT 52.000 126.900 52.900 127.100 ;
        RECT 52.100 126.800 52.900 126.900 ;
        RECT 47.800 126.100 48.200 126.200 ;
        RECT 45.400 125.800 46.200 126.100 ;
        RECT 47.000 125.800 48.200 126.100 ;
        RECT 51.000 125.800 51.800 126.200 ;
        RECT 45.800 125.600 46.200 125.800 ;
        RECT 44.600 125.100 45.000 125.200 ;
        RECT 47.800 125.100 48.100 125.800 ;
        RECT 43.500 124.800 44.000 125.100 ;
        RECT 44.300 124.800 45.000 125.100 ;
        RECT 45.400 124.800 47.400 125.100 ;
        RECT 30.500 121.100 30.900 124.700 ;
        RECT 32.700 124.400 34.500 124.700 ;
        RECT 32.700 124.100 33.000 124.400 ;
        RECT 32.600 121.100 33.000 124.100 ;
        RECT 34.200 124.100 34.500 124.400 ;
        RECT 35.100 124.500 36.900 124.600 ;
        RECT 37.400 124.500 37.700 124.800 ;
        RECT 35.100 124.300 37.000 124.500 ;
        RECT 35.100 124.100 35.400 124.300 ;
        RECT 34.200 121.400 34.600 124.100 ;
        RECT 35.000 121.700 35.400 124.100 ;
        RECT 35.800 121.400 36.200 124.000 ;
        RECT 36.600 121.500 37.000 124.300 ;
        RECT 37.400 121.700 37.800 124.500 ;
        RECT 34.200 121.100 36.200 121.400 ;
        RECT 36.700 121.400 37.000 121.500 ;
        RECT 38.200 121.500 38.600 124.500 ;
        RECT 39.100 123.500 39.400 124.800 ;
        RECT 39.800 124.100 40.200 124.600 ;
        RECT 40.600 124.100 41.000 124.200 ;
        RECT 39.800 123.800 41.000 124.100 ;
        RECT 39.100 123.200 40.900 123.500 ;
        RECT 39.100 123.100 39.400 123.200 ;
        RECT 38.200 121.400 38.500 121.500 ;
        RECT 36.700 121.100 38.500 121.400 ;
        RECT 39.000 121.100 39.400 123.100 ;
        RECT 40.600 123.100 40.900 123.200 ;
        RECT 40.600 121.100 41.000 123.100 ;
        RECT 43.500 121.100 43.900 124.800 ;
        RECT 44.300 124.200 44.600 124.800 ;
        RECT 44.200 123.800 44.600 124.200 ;
        RECT 45.400 121.100 45.800 124.800 ;
        RECT 47.000 121.100 47.400 124.800 ;
        RECT 47.800 121.100 48.200 125.100 ;
        RECT 50.200 124.800 50.600 125.600 ;
        RECT 52.600 125.200 52.900 126.800 ;
        RECT 53.500 126.900 54.400 127.100 ;
        RECT 53.500 126.800 54.300 126.900 ;
        RECT 53.500 125.200 53.800 126.800 ;
        RECT 54.600 125.800 55.400 126.200 ;
        RECT 52.600 124.800 53.000 125.200 ;
        RECT 53.400 124.800 53.800 125.200 ;
        RECT 55.800 124.800 56.200 125.600 ;
        RECT 58.800 125.200 59.100 127.800 ;
        RECT 63.100 127.700 64.900 127.900 ;
        RECT 63.400 127.200 63.800 127.400 ;
        RECT 65.400 127.200 65.700 127.900 ;
        RECT 66.200 127.800 66.600 128.600 ;
        RECT 60.200 127.100 61.000 127.200 ;
        RECT 60.200 126.800 62.500 127.100 ;
        RECT 63.000 126.900 63.800 127.200 ;
        RECT 63.000 126.800 63.400 126.900 ;
        RECT 64.500 126.800 65.800 127.200 ;
        RECT 66.200 127.100 66.600 127.200 ;
        RECT 67.000 127.100 67.400 129.900 ;
        RECT 66.200 126.800 67.400 127.100 ;
        RECT 69.600 127.100 70.000 129.900 ;
        RECT 69.600 126.900 70.500 127.100 ;
        RECT 69.700 126.800 70.500 126.900 ;
        RECT 62.200 126.200 62.500 126.800 ;
        RECT 59.400 125.800 60.200 126.200 ;
        RECT 62.200 126.100 62.600 126.200 ;
        RECT 63.800 126.100 64.200 126.600 ;
        RECT 62.200 125.800 64.200 126.100 ;
        RECT 57.400 124.900 59.100 125.200 ;
        RECT 64.500 125.100 64.800 126.800 ;
        RECT 65.400 125.100 65.800 125.200 ;
        RECT 57.400 124.800 57.800 124.900 ;
        RECT 51.800 123.800 52.200 124.600 ;
        RECT 52.600 124.200 52.900 124.800 ;
        RECT 52.600 123.800 53.000 124.200 ;
        RECT 52.600 123.500 52.900 123.800 ;
        RECT 51.100 123.200 52.900 123.500 ;
        RECT 51.100 123.100 51.400 123.200 ;
        RECT 51.000 121.100 51.400 123.100 ;
        RECT 52.600 123.100 52.900 123.200 ;
        RECT 53.500 123.500 53.800 124.800 ;
        RECT 54.200 123.800 54.600 124.600 ;
        RECT 57.500 124.500 57.800 124.800 ;
        RECT 64.300 124.800 64.800 125.100 ;
        RECT 65.100 124.800 65.800 125.100 ;
        RECT 58.300 124.500 60.100 124.600 ;
        RECT 53.500 123.200 55.300 123.500 ;
        RECT 53.500 123.100 53.800 123.200 ;
        RECT 52.600 121.100 53.000 123.100 ;
        RECT 53.400 121.100 53.800 123.100 ;
        RECT 55.000 123.100 55.300 123.200 ;
        RECT 55.000 121.100 55.400 123.100 ;
        RECT 56.600 121.500 57.000 124.500 ;
        RECT 57.400 121.700 57.800 124.500 ;
        RECT 58.200 124.300 60.100 124.500 ;
        RECT 56.700 121.400 57.000 121.500 ;
        RECT 58.200 121.500 58.600 124.300 ;
        RECT 59.800 124.100 60.100 124.300 ;
        RECT 60.700 124.400 62.500 124.700 ;
        RECT 60.700 124.100 61.000 124.400 ;
        RECT 58.200 121.400 58.500 121.500 ;
        RECT 56.700 121.100 58.500 121.400 ;
        RECT 59.000 121.400 59.400 124.000 ;
        RECT 59.800 121.700 60.200 124.100 ;
        RECT 60.600 121.400 61.000 124.100 ;
        RECT 59.000 121.100 61.000 121.400 ;
        RECT 62.200 124.100 62.500 124.400 ;
        RECT 62.200 121.100 62.600 124.100 ;
        RECT 64.300 121.100 64.700 124.800 ;
        RECT 65.100 124.200 65.400 124.800 ;
        RECT 65.000 123.800 65.400 124.200 ;
        RECT 67.000 121.100 67.400 126.800 ;
        RECT 68.600 125.800 69.400 126.200 ;
        RECT 67.800 124.800 68.200 125.600 ;
        RECT 70.200 125.200 70.500 126.800 ;
        RECT 70.200 124.800 70.600 125.200 ;
        RECT 69.400 123.800 69.800 124.600 ;
        RECT 70.200 124.200 70.500 124.800 ;
        RECT 70.200 123.800 70.600 124.200 ;
        RECT 70.200 123.500 70.500 123.800 ;
        RECT 68.700 123.200 70.500 123.500 ;
        RECT 68.700 123.100 69.000 123.200 ;
        RECT 68.600 121.100 69.000 123.100 ;
        RECT 70.200 123.100 70.500 123.200 ;
        RECT 70.200 121.100 70.600 123.100 ;
        RECT 71.000 121.100 71.400 129.900 ;
        RECT 71.800 127.800 72.200 128.600 ;
        RECT 73.200 127.100 73.600 129.900 ;
        RECT 72.700 126.900 73.600 127.100 ;
        RECT 76.600 127.600 77.000 129.900 ;
        RECT 78.200 127.600 78.600 129.900 ;
        RECT 76.600 127.200 78.600 127.600 ;
        RECT 72.700 126.800 73.500 126.900 ;
        RECT 72.700 125.200 73.000 126.800 ;
        RECT 73.800 125.800 74.600 126.200 ;
        RECT 76.600 125.800 77.000 127.200 ;
        RECT 78.200 126.800 78.600 127.200 ;
        RECT 80.400 127.100 80.800 129.900 ;
        RECT 79.900 126.900 80.800 127.100 ;
        RECT 83.000 126.900 83.400 129.900 ;
        RECT 86.200 128.300 86.600 129.900 ;
        RECT 87.000 128.500 87.400 129.900 ;
        RECT 87.800 128.500 88.200 129.900 ;
        RECT 88.600 128.500 89.000 129.900 ;
        RECT 90.200 128.500 90.600 129.900 ;
        RECT 91.800 128.500 92.200 129.900 ;
        RECT 92.600 128.500 93.000 129.900 ;
        RECT 93.400 128.500 93.800 129.900 ;
        RECT 94.200 128.500 94.600 129.900 ;
        RECT 85.300 127.900 86.600 128.300 ;
        RECT 95.000 128.300 95.400 129.900 ;
        RECT 88.300 127.900 90.600 128.200 ;
        RECT 85.300 127.600 85.700 127.900 ;
        RECT 84.200 127.200 85.700 127.600 ;
        RECT 79.900 126.800 80.700 126.900 ;
        RECT 72.600 124.800 73.000 125.200 ;
        RECT 74.200 125.100 74.600 125.200 ;
        RECT 75.000 125.100 75.400 125.600 ;
        RECT 74.200 124.800 75.400 125.100 ;
        RECT 76.600 125.400 78.600 125.800 ;
        RECT 72.700 123.500 73.000 124.800 ;
        RECT 73.400 123.800 73.800 124.600 ;
        RECT 72.700 123.200 74.500 123.500 ;
        RECT 72.700 123.100 73.000 123.200 ;
        RECT 72.600 121.100 73.000 123.100 ;
        RECT 74.200 123.100 74.500 123.200 ;
        RECT 74.200 121.100 74.600 123.100 ;
        RECT 76.600 121.100 77.000 125.400 ;
        RECT 78.200 121.100 78.600 125.400 ;
        RECT 79.900 125.200 80.200 126.800 ;
        RECT 83.000 126.500 87.400 126.900 ;
        RECT 88.300 126.700 88.700 127.900 ;
        RECT 90.200 127.800 90.600 127.900 ;
        RECT 93.300 127.800 93.800 128.200 ;
        RECT 95.000 127.900 96.200 128.300 ;
        RECT 89.400 126.800 89.800 127.600 ;
        RECT 90.200 127.400 90.600 127.500 ;
        RECT 90.200 127.100 92.400 127.400 ;
        RECT 92.000 127.000 92.400 127.100 ;
        RECT 81.000 125.800 81.800 126.200 ;
        RECT 79.800 124.800 80.200 125.200 ;
        RECT 82.200 124.800 82.600 125.600 ;
        RECT 79.900 123.500 80.200 124.800 ;
        RECT 80.600 123.800 81.000 124.600 ;
        RECT 83.000 123.700 83.400 126.500 ;
        RECT 87.700 126.300 88.700 126.700 ;
        RECT 90.600 126.300 92.200 126.700 ;
        RECT 93.400 126.400 93.800 127.800 ;
        RECT 95.800 127.600 96.200 127.900 ;
        RECT 95.800 127.300 96.700 127.600 ;
        RECT 95.000 126.800 95.400 127.200 ;
        RECT 95.000 126.300 95.300 126.800 ;
        RECT 96.300 126.700 96.700 127.300 ;
        RECT 98.200 127.300 98.600 129.900 ;
        RECT 99.000 128.000 99.400 129.900 ;
        RECT 99.000 127.600 99.500 128.000 ;
        RECT 98.200 127.000 98.800 127.300 ;
        RECT 96.300 126.300 98.200 126.700 ;
        RECT 83.700 126.000 84.100 126.100 ;
        RECT 84.600 126.000 85.000 126.200 ;
        RECT 86.200 126.000 86.600 126.200 ;
        RECT 95.000 126.000 95.400 126.300 ;
        RECT 98.500 126.000 98.800 127.000 ;
        RECT 83.700 125.700 95.400 126.000 ;
        RECT 98.400 125.700 98.800 126.000 ;
        RECT 98.400 124.800 98.700 125.700 ;
        RECT 99.100 125.400 99.500 127.600 ;
        RECT 87.800 124.700 88.200 124.800 ;
        RECT 85.500 124.500 88.200 124.700 ;
        RECT 85.100 124.400 88.200 124.500 ;
        RECT 88.700 124.500 93.000 124.800 ;
        RECT 83.800 124.000 84.600 124.400 ;
        RECT 85.100 124.100 85.800 124.400 ;
        RECT 88.700 124.100 89.000 124.500 ;
        RECT 92.600 124.400 93.000 124.500 ;
        RECT 94.200 124.500 98.700 124.800 ;
        RECT 94.200 124.400 94.600 124.500 ;
        RECT 84.300 123.800 84.600 124.000 ;
        RECT 86.100 123.800 89.000 124.100 ;
        RECT 89.300 123.800 90.600 124.200 ;
        RECT 79.900 123.200 81.700 123.500 ;
        RECT 83.000 123.400 84.000 123.700 ;
        RECT 84.300 123.400 86.400 123.800 ;
        RECT 79.900 123.100 80.200 123.200 ;
        RECT 79.800 121.100 80.200 123.100 ;
        RECT 81.400 123.100 81.700 123.200 ;
        RECT 83.700 123.100 84.000 123.400 ;
        RECT 81.400 121.100 81.800 123.100 ;
        RECT 83.700 122.800 84.200 123.100 ;
        RECT 83.800 121.100 84.200 122.800 ;
        RECT 85.400 121.100 85.800 123.400 ;
        RECT 87.000 121.100 87.400 122.500 ;
        RECT 87.800 121.100 88.200 122.500 ;
        RECT 88.600 121.100 89.000 123.500 ;
        RECT 90.200 121.100 90.600 123.500 ;
        RECT 91.800 121.100 92.200 124.200 ;
        RECT 95.800 123.800 97.100 124.200 ;
        RECT 93.400 123.400 95.500 123.800 ;
        RECT 92.600 121.100 93.000 122.500 ;
        RECT 93.400 121.100 93.800 122.500 ;
        RECT 94.200 121.100 94.600 122.500 ;
        RECT 95.800 121.100 96.200 123.800 ;
        RECT 98.400 123.700 98.700 124.500 ;
        RECT 97.400 123.400 98.700 123.700 ;
        RECT 99.000 125.000 99.500 125.400 ;
        RECT 102.200 126.900 102.600 129.900 ;
        RECT 105.400 128.300 105.800 129.900 ;
        RECT 106.200 128.500 106.600 129.900 ;
        RECT 107.000 128.500 107.400 129.900 ;
        RECT 107.800 128.500 108.200 129.900 ;
        RECT 109.400 128.500 109.800 129.900 ;
        RECT 111.000 128.500 111.400 129.900 ;
        RECT 111.800 128.500 112.200 129.900 ;
        RECT 112.600 128.500 113.000 129.900 ;
        RECT 113.400 128.500 113.800 129.900 ;
        RECT 104.500 127.900 105.800 128.300 ;
        RECT 114.200 128.300 114.600 129.900 ;
        RECT 107.500 127.900 109.800 128.200 ;
        RECT 104.500 127.600 104.900 127.900 ;
        RECT 103.400 127.200 104.900 127.600 ;
        RECT 102.200 126.500 106.600 126.900 ;
        RECT 107.500 126.700 107.900 127.900 ;
        RECT 109.400 127.800 109.800 127.900 ;
        RECT 112.500 127.800 113.000 128.200 ;
        RECT 114.200 127.900 115.400 128.300 ;
        RECT 108.600 126.800 109.000 127.600 ;
        RECT 109.400 127.400 109.800 127.500 ;
        RECT 109.400 127.100 111.600 127.400 ;
        RECT 111.200 127.000 111.600 127.100 ;
        RECT 97.400 121.100 97.800 123.400 ;
        RECT 99.000 121.100 99.400 125.000 ;
        RECT 102.200 123.700 102.600 126.500 ;
        RECT 106.900 126.300 107.900 126.700 ;
        RECT 109.800 126.300 111.400 126.700 ;
        RECT 112.600 126.400 113.000 127.800 ;
        RECT 115.000 127.600 115.400 127.900 ;
        RECT 115.000 127.300 115.900 127.600 ;
        RECT 115.500 126.700 115.900 127.300 ;
        RECT 117.400 127.300 117.800 129.900 ;
        RECT 118.200 128.000 118.600 129.900 ;
        RECT 118.200 127.600 118.700 128.000 ;
        RECT 117.400 127.000 118.000 127.300 ;
        RECT 115.500 126.300 117.400 126.700 ;
        RECT 102.900 126.000 103.300 126.100 ;
        RECT 103.800 126.000 104.200 126.200 ;
        RECT 105.400 126.000 105.800 126.200 ;
        RECT 114.200 126.000 114.600 126.300 ;
        RECT 117.700 126.000 118.000 127.000 ;
        RECT 102.900 125.700 114.600 126.000 ;
        RECT 117.600 125.700 118.000 126.000 ;
        RECT 117.600 124.800 117.900 125.700 ;
        RECT 118.300 125.400 118.700 127.600 ;
        RECT 107.000 124.700 107.400 124.800 ;
        RECT 104.700 124.500 107.400 124.700 ;
        RECT 104.300 124.400 107.400 124.500 ;
        RECT 107.900 124.500 112.200 124.800 ;
        RECT 103.000 124.000 103.800 124.400 ;
        RECT 104.300 124.100 105.000 124.400 ;
        RECT 107.900 124.100 108.200 124.500 ;
        RECT 111.800 124.400 112.200 124.500 ;
        RECT 113.400 124.500 117.900 124.800 ;
        RECT 113.400 124.400 113.800 124.500 ;
        RECT 103.500 123.800 103.800 124.000 ;
        RECT 105.300 123.800 108.200 124.100 ;
        RECT 108.500 123.800 109.800 124.200 ;
        RECT 102.200 123.400 103.200 123.700 ;
        RECT 103.500 123.400 105.600 123.800 ;
        RECT 102.900 123.100 103.200 123.400 ;
        RECT 102.900 122.800 103.400 123.100 ;
        RECT 103.000 121.100 103.400 122.800 ;
        RECT 104.600 121.100 105.000 123.400 ;
        RECT 106.200 121.100 106.600 122.500 ;
        RECT 107.000 121.100 107.400 122.500 ;
        RECT 107.800 121.100 108.200 123.500 ;
        RECT 109.400 121.100 109.800 123.500 ;
        RECT 111.000 121.100 111.400 124.200 ;
        RECT 115.000 123.800 116.300 124.200 ;
        RECT 112.600 123.400 114.700 123.800 ;
        RECT 111.800 121.100 112.200 122.500 ;
        RECT 112.600 121.100 113.000 122.500 ;
        RECT 113.400 121.100 113.800 122.500 ;
        RECT 115.000 121.100 115.400 123.800 ;
        RECT 117.600 123.700 117.900 124.500 ;
        RECT 116.600 123.400 117.900 123.700 ;
        RECT 118.200 125.000 118.700 125.400 ;
        RECT 116.600 121.100 117.000 123.400 ;
        RECT 118.200 121.100 118.600 125.000 ;
        RECT 119.800 121.100 120.200 129.900 ;
        RECT 120.600 127.800 121.000 128.600 ;
        RECT 121.400 126.900 121.800 129.900 ;
        RECT 124.600 128.300 125.000 129.900 ;
        RECT 125.400 128.500 125.800 129.900 ;
        RECT 126.200 128.500 126.600 129.900 ;
        RECT 127.000 128.500 127.400 129.900 ;
        RECT 128.600 128.500 129.000 129.900 ;
        RECT 130.200 128.500 130.600 129.900 ;
        RECT 131.000 128.500 131.400 129.900 ;
        RECT 131.800 128.500 132.200 129.900 ;
        RECT 132.600 128.500 133.000 129.900 ;
        RECT 123.700 127.900 125.000 128.300 ;
        RECT 133.400 128.300 133.800 129.900 ;
        RECT 126.700 127.900 129.000 128.200 ;
        RECT 123.700 127.600 124.100 127.900 ;
        RECT 122.600 127.200 124.100 127.600 ;
        RECT 121.400 126.500 125.800 126.900 ;
        RECT 126.700 126.700 127.100 127.900 ;
        RECT 128.600 127.800 129.000 127.900 ;
        RECT 131.700 127.800 132.200 128.200 ;
        RECT 133.400 127.900 134.600 128.300 ;
        RECT 127.800 126.800 128.200 127.600 ;
        RECT 128.600 127.400 129.000 127.500 ;
        RECT 128.600 127.100 130.800 127.400 ;
        RECT 130.400 127.000 130.800 127.100 ;
        RECT 121.400 123.700 121.800 126.500 ;
        RECT 126.100 126.300 127.100 126.700 ;
        RECT 129.000 126.300 130.600 126.700 ;
        RECT 131.800 126.400 132.200 127.800 ;
        RECT 134.200 127.600 134.600 127.900 ;
        RECT 134.200 127.300 135.100 127.600 ;
        RECT 134.700 126.700 135.100 127.300 ;
        RECT 136.600 127.300 137.000 129.900 ;
        RECT 137.400 128.100 137.800 129.900 ;
        RECT 138.200 128.100 138.600 128.200 ;
        RECT 137.400 127.800 138.600 128.100 ;
        RECT 137.400 127.600 137.900 127.800 ;
        RECT 136.600 127.000 137.200 127.300 ;
        RECT 134.700 126.300 136.600 126.700 ;
        RECT 122.100 126.000 122.500 126.100 ;
        RECT 123.000 126.000 123.400 126.200 ;
        RECT 124.600 126.000 125.000 126.200 ;
        RECT 133.400 126.000 133.800 126.300 ;
        RECT 136.900 126.000 137.200 127.000 ;
        RECT 122.100 125.700 133.800 126.000 ;
        RECT 136.800 125.700 137.200 126.000 ;
        RECT 137.500 126.100 137.900 127.600 ;
        RECT 139.000 127.600 139.400 129.900 ;
        RECT 141.400 127.600 141.800 129.900 ;
        RECT 143.800 127.600 144.200 129.900 ;
        RECT 139.000 127.300 140.100 127.600 ;
        RECT 141.400 127.300 142.500 127.600 ;
        RECT 143.800 127.300 144.900 127.600 ;
        RECT 139.000 126.100 139.400 126.600 ;
        RECT 137.500 125.800 139.400 126.100 ;
        RECT 139.800 125.800 140.100 127.300 ;
        RECT 141.400 125.800 141.800 126.600 ;
        RECT 142.200 125.800 142.500 127.300 ;
        RECT 143.800 125.800 144.200 126.600 ;
        RECT 144.600 125.800 144.900 127.300 ;
        RECT 136.800 124.800 137.100 125.700 ;
        RECT 137.500 125.400 137.900 125.800 ;
        RECT 126.200 124.700 126.600 124.800 ;
        RECT 123.900 124.500 126.600 124.700 ;
        RECT 123.500 124.400 126.600 124.500 ;
        RECT 127.100 124.500 131.400 124.800 ;
        RECT 122.200 124.000 123.000 124.400 ;
        RECT 123.500 124.100 124.200 124.400 ;
        RECT 127.100 124.100 127.400 124.500 ;
        RECT 131.000 124.400 131.400 124.500 ;
        RECT 132.600 124.500 137.100 124.800 ;
        RECT 132.600 124.400 133.000 124.500 ;
        RECT 122.700 123.800 123.000 124.000 ;
        RECT 124.500 123.800 127.400 124.100 ;
        RECT 127.700 123.800 129.000 124.200 ;
        RECT 121.400 123.400 122.400 123.700 ;
        RECT 122.700 123.400 124.800 123.800 ;
        RECT 122.100 123.100 122.400 123.400 ;
        RECT 122.100 122.800 122.600 123.100 ;
        RECT 122.200 121.100 122.600 122.800 ;
        RECT 123.800 121.100 124.200 123.400 ;
        RECT 125.400 121.100 125.800 122.500 ;
        RECT 126.200 121.100 126.600 122.500 ;
        RECT 127.000 121.100 127.400 123.500 ;
        RECT 128.600 121.100 129.000 123.500 ;
        RECT 130.200 121.100 130.600 124.200 ;
        RECT 134.200 123.800 135.500 124.200 ;
        RECT 131.800 123.400 133.900 123.800 ;
        RECT 131.000 121.100 131.400 122.500 ;
        RECT 131.800 121.100 132.200 122.500 ;
        RECT 132.600 121.100 133.000 122.500 ;
        RECT 134.200 121.100 134.600 123.800 ;
        RECT 136.800 123.700 137.100 124.500 ;
        RECT 135.800 123.400 137.100 123.700 ;
        RECT 137.400 125.000 137.900 125.400 ;
        RECT 139.800 125.400 140.400 125.800 ;
        RECT 142.200 125.400 142.800 125.800 ;
        RECT 144.600 125.400 145.200 125.800 ;
        RECT 139.800 125.100 140.100 125.400 ;
        RECT 142.200 125.100 142.500 125.400 ;
        RECT 144.600 125.100 144.900 125.400 ;
        RECT 135.800 121.100 136.200 123.400 ;
        RECT 137.400 121.100 137.800 125.000 ;
        RECT 139.000 124.800 140.100 125.100 ;
        RECT 141.400 124.800 142.500 125.100 ;
        RECT 143.800 124.800 144.900 125.100 ;
        RECT 139.000 121.100 139.400 124.800 ;
        RECT 141.400 121.100 141.800 124.800 ;
        RECT 143.800 121.100 144.200 124.800 ;
        RECT 147.000 121.100 147.400 129.900 ;
        RECT 148.100 128.200 148.500 129.900 ;
        RECT 148.100 127.900 149.000 128.200 ;
        RECT 147.800 124.400 148.200 125.200 ;
        RECT 148.600 121.100 149.000 127.900 ;
        RECT 0.600 117.900 1.000 119.900 ;
        RECT 0.700 117.800 1.000 117.900 ;
        RECT 2.200 117.900 2.600 119.900 ;
        RECT 3.800 117.900 4.200 119.900 ;
        RECT 2.200 117.800 2.500 117.900 ;
        RECT 0.700 117.500 2.500 117.800 ;
        RECT 3.900 117.800 4.200 117.900 ;
        RECT 5.400 117.900 5.800 119.900 ;
        RECT 5.400 117.800 5.700 117.900 ;
        RECT 3.900 117.500 5.700 117.800 ;
        RECT 0.700 116.200 1.000 117.500 ;
        RECT 1.400 116.400 1.800 117.200 ;
        RECT 3.900 116.200 4.200 117.500 ;
        RECT 4.600 116.400 5.000 117.200 ;
        RECT 7.300 116.300 7.700 119.900 ;
        RECT 9.400 117.900 9.800 119.900 ;
        RECT 9.500 117.800 9.800 117.900 ;
        RECT 11.000 117.900 11.400 119.900 ;
        RECT 11.000 117.800 11.300 117.900 ;
        RECT 9.500 117.500 11.300 117.800 ;
        RECT 0.600 115.800 1.000 116.200 ;
        RECT 0.700 114.200 1.000 115.800 ;
        RECT 3.000 115.400 3.400 116.200 ;
        RECT 3.800 115.800 4.200 116.200 ;
        RECT 3.900 115.200 4.200 115.800 ;
        RECT 6.200 115.400 6.600 116.200 ;
        RECT 7.300 115.900 8.200 116.300 ;
        RECT 9.500 116.200 9.800 117.500 ;
        RECT 1.800 114.800 2.600 115.200 ;
        RECT 3.800 114.800 4.200 115.200 ;
        RECT 5.000 114.800 5.800 115.200 ;
        RECT 7.000 114.800 7.400 115.600 ;
        RECT 3.900 114.200 4.200 114.800 ;
        RECT 7.000 114.200 7.300 114.800 ;
        RECT 7.800 114.200 8.100 115.900 ;
        RECT 9.400 115.800 9.800 116.200 ;
        RECT 10.200 117.100 10.600 117.200 ;
        RECT 12.600 117.100 13.000 117.200 ;
        RECT 10.200 116.800 13.000 117.100 ;
        RECT 10.200 115.800 10.600 116.800 ;
        RECT 9.500 114.200 9.800 115.800 ;
        RECT 11.800 115.400 12.200 116.200 ;
        RECT 12.600 115.800 13.000 116.800 ;
        RECT 10.600 114.800 11.400 115.200 ;
        RECT 0.700 114.100 1.500 114.200 ;
        RECT 3.900 114.100 4.700 114.200 ;
        RECT 0.700 113.900 1.600 114.100 ;
        RECT 3.900 113.900 4.800 114.100 ;
        RECT 1.200 111.100 1.600 113.900 ;
        RECT 4.400 111.100 4.800 113.900 ;
        RECT 7.000 113.800 7.400 114.200 ;
        RECT 7.800 113.800 8.200 114.200 ;
        RECT 9.500 114.100 10.300 114.200 ;
        RECT 9.500 113.900 10.400 114.100 ;
        RECT 7.800 112.200 8.100 113.800 ;
        RECT 8.600 112.400 9.000 113.200 ;
        RECT 7.800 111.100 8.200 112.200 ;
        RECT 10.000 111.100 10.400 113.900 ;
        RECT 13.400 113.100 13.800 119.900 ;
        RECT 15.800 117.900 16.200 119.900 ;
        RECT 15.900 117.800 16.200 117.900 ;
        RECT 17.400 117.900 17.800 119.900 ;
        RECT 17.400 117.800 17.700 117.900 ;
        RECT 15.900 117.500 17.700 117.800 ;
        RECT 15.800 117.100 16.200 117.200 ;
        RECT 16.600 117.100 17.000 117.200 ;
        RECT 15.800 116.800 17.000 117.100 ;
        RECT 16.600 116.400 17.000 116.800 ;
        RECT 17.400 116.200 17.700 117.500 ;
        RECT 18.600 116.800 19.000 117.200 ;
        RECT 18.600 116.200 18.900 116.800 ;
        RECT 19.300 116.200 19.700 119.900 ;
        RECT 14.200 116.100 14.600 116.200 ;
        RECT 15.000 116.100 15.400 116.200 ;
        RECT 14.200 115.800 15.400 116.100 ;
        RECT 15.000 115.400 15.400 115.800 ;
        RECT 17.400 115.800 17.800 116.200 ;
        RECT 18.200 115.900 18.900 116.200 ;
        RECT 19.200 115.900 19.700 116.200 ;
        RECT 18.200 115.800 18.600 115.900 ;
        RECT 15.800 114.800 17.000 115.200 ;
        RECT 17.400 114.200 17.700 115.800 ;
        RECT 19.200 114.200 19.500 115.900 ;
        RECT 19.800 115.100 20.200 115.200 ;
        RECT 21.400 115.100 21.800 119.900 ;
        RECT 23.000 116.200 23.400 119.900 ;
        RECT 24.600 116.200 25.000 119.900 ;
        RECT 23.000 115.900 25.000 116.200 ;
        RECT 25.400 115.900 25.800 119.900 ;
        RECT 27.500 117.200 27.900 119.900 ;
        RECT 27.000 116.800 27.900 117.200 ;
        RECT 28.200 116.800 28.600 117.200 ;
        RECT 27.500 116.200 27.900 116.800 ;
        RECT 28.300 116.200 28.600 116.800 ;
        RECT 29.400 116.200 29.800 119.900 ;
        RECT 31.000 116.200 31.400 119.900 ;
        RECT 27.500 115.900 28.000 116.200 ;
        RECT 28.300 115.900 29.000 116.200 ;
        RECT 29.400 115.900 31.400 116.200 ;
        RECT 31.800 115.900 32.200 119.900 ;
        RECT 32.600 117.900 33.000 119.900 ;
        RECT 32.700 117.800 33.000 117.900 ;
        RECT 34.200 117.900 34.600 119.900 ;
        RECT 36.600 117.900 37.000 119.900 ;
        RECT 34.200 117.800 34.500 117.900 ;
        RECT 32.700 117.500 34.500 117.800 ;
        RECT 36.700 117.800 37.000 117.900 ;
        RECT 38.200 117.900 38.600 119.900 ;
        RECT 40.100 119.200 40.500 119.900 ;
        RECT 40.100 118.800 41.000 119.200 ;
        RECT 38.200 117.800 38.500 117.900 ;
        RECT 36.700 117.500 38.500 117.800 ;
        RECT 32.700 116.200 33.000 117.500 ;
        RECT 33.400 116.400 33.800 117.200 ;
        RECT 37.400 116.400 37.800 117.200 ;
        RECT 38.200 116.200 38.500 117.500 ;
        RECT 39.400 116.800 39.800 117.200 ;
        RECT 39.400 116.200 39.700 116.800 ;
        RECT 40.100 116.200 40.500 118.800 ;
        RECT 43.000 117.900 43.400 119.900 ;
        RECT 43.100 117.800 43.400 117.900 ;
        RECT 44.600 117.900 45.000 119.900 ;
        RECT 44.600 117.800 44.900 117.900 ;
        RECT 43.100 117.500 44.900 117.800 ;
        RECT 43.800 116.400 44.200 117.200 ;
        RECT 44.600 116.200 44.900 117.500 ;
        RECT 23.400 115.200 23.800 115.400 ;
        RECT 25.400 115.200 25.700 115.900 ;
        RECT 19.800 114.800 21.800 115.100 ;
        RECT 23.000 114.900 23.800 115.200 ;
        RECT 24.600 114.900 25.800 115.200 ;
        RECT 23.000 114.800 23.400 114.900 ;
        RECT 19.800 114.400 20.200 114.800 ;
        RECT 14.200 113.400 14.600 114.200 ;
        RECT 16.900 114.100 17.700 114.200 ;
        RECT 16.800 113.900 17.700 114.100 ;
        RECT 12.900 112.800 13.800 113.100 ;
        RECT 12.900 112.200 13.300 112.800 ;
        RECT 12.600 111.800 13.300 112.200 ;
        RECT 12.900 111.100 13.300 111.800 ;
        RECT 16.800 111.100 17.200 113.900 ;
        RECT 18.200 113.800 19.500 114.200 ;
        RECT 20.600 114.100 21.000 114.200 ;
        RECT 20.200 113.800 21.000 114.100 ;
        RECT 18.300 113.200 18.600 113.800 ;
        RECT 20.200 113.600 20.600 113.800 ;
        RECT 18.200 111.100 18.600 113.200 ;
        RECT 19.100 113.100 20.900 113.300 ;
        RECT 19.000 113.000 21.000 113.100 ;
        RECT 19.000 111.100 19.400 113.000 ;
        RECT 20.600 111.100 21.000 113.000 ;
        RECT 21.400 111.100 21.800 114.800 ;
        RECT 22.200 114.100 22.600 114.200 ;
        RECT 23.000 114.100 23.400 114.200 ;
        RECT 22.200 113.800 23.400 114.100 ;
        RECT 23.800 113.800 24.200 114.600 ;
        RECT 22.200 113.400 22.600 113.800 ;
        RECT 24.600 113.100 24.900 114.900 ;
        RECT 25.400 114.800 25.800 114.900 ;
        RECT 26.200 115.100 26.600 115.200 ;
        RECT 27.000 115.100 27.400 115.200 ;
        RECT 26.200 114.800 27.400 115.100 ;
        RECT 27.000 114.400 27.400 114.800 ;
        RECT 27.700 114.200 28.000 115.900 ;
        RECT 28.600 115.800 29.000 115.900 ;
        RECT 29.800 115.200 30.200 115.400 ;
        RECT 31.800 115.200 32.100 115.900 ;
        RECT 32.600 115.800 33.000 116.200 ;
        RECT 29.400 114.900 30.200 115.200 ;
        RECT 31.000 114.900 32.200 115.200 ;
        RECT 29.400 114.800 29.800 114.900 ;
        RECT 26.200 114.100 26.600 114.200 ;
        RECT 26.200 113.800 27.000 114.100 ;
        RECT 27.700 113.800 29.000 114.200 ;
        RECT 30.200 113.800 30.600 114.600 ;
        RECT 26.600 113.600 27.000 113.800 ;
        RECT 24.600 111.100 25.000 113.100 ;
        RECT 25.400 112.800 25.800 113.200 ;
        RECT 26.300 113.100 28.100 113.300 ;
        RECT 28.600 113.100 28.900 113.800 ;
        RECT 31.000 113.100 31.300 114.900 ;
        RECT 31.800 114.800 32.200 114.900 ;
        RECT 32.700 114.200 33.000 115.800 ;
        RECT 35.000 115.400 35.400 116.200 ;
        RECT 35.800 115.400 36.200 116.200 ;
        RECT 38.200 115.800 38.600 116.200 ;
        RECT 39.000 115.900 39.700 116.200 ;
        RECT 40.000 115.900 40.500 116.200 ;
        RECT 39.000 115.800 39.400 115.900 ;
        RECT 33.800 114.800 34.600 115.200 ;
        RECT 36.600 114.800 37.400 115.200 ;
        RECT 38.200 114.200 38.500 115.800 ;
        RECT 40.000 114.200 40.300 115.900 ;
        RECT 42.200 115.400 42.600 116.200 ;
        RECT 44.600 115.800 45.000 116.200 ;
        RECT 45.400 115.900 45.800 119.900 ;
        RECT 46.200 116.200 46.600 119.900 ;
        RECT 47.800 116.200 48.200 119.900 ;
        RECT 46.200 115.900 48.200 116.200 ;
        RECT 40.600 114.400 41.000 115.200 ;
        RECT 43.000 114.800 43.800 115.200 ;
        RECT 44.600 114.200 44.900 115.800 ;
        RECT 45.500 115.200 45.800 115.900 ;
        RECT 47.400 115.200 47.800 115.400 ;
        RECT 45.400 114.900 46.600 115.200 ;
        RECT 47.400 115.100 48.200 115.200 ;
        RECT 50.200 115.100 50.600 119.900 ;
        RECT 47.400 114.900 50.600 115.100 ;
        RECT 45.400 114.800 45.800 114.900 ;
        RECT 32.700 113.900 33.800 114.200 ;
        RECT 37.700 114.100 38.500 114.200 ;
        RECT 33.200 113.800 33.800 113.900 ;
        RECT 37.600 113.900 38.500 114.100 ;
        RECT 26.200 113.000 28.200 113.100 ;
        RECT 25.300 112.400 25.700 112.800 ;
        RECT 26.200 111.100 26.600 113.000 ;
        RECT 27.800 111.100 28.200 113.000 ;
        RECT 28.600 111.100 29.000 113.100 ;
        RECT 31.000 111.100 31.400 113.100 ;
        RECT 31.800 112.800 32.200 113.200 ;
        RECT 31.700 112.400 32.100 112.800 ;
        RECT 33.200 111.100 33.600 113.800 ;
        RECT 37.600 111.100 38.000 113.900 ;
        RECT 39.000 113.800 40.300 114.200 ;
        RECT 41.400 114.100 41.800 114.200 ;
        RECT 44.100 114.100 44.900 114.200 ;
        RECT 41.000 113.800 41.800 114.100 ;
        RECT 44.000 113.900 44.900 114.100 ;
        RECT 39.100 113.100 39.400 113.800 ;
        RECT 41.000 113.600 41.400 113.800 ;
        RECT 39.900 113.100 41.700 113.300 ;
        RECT 39.000 111.100 39.400 113.100 ;
        RECT 39.800 113.000 41.800 113.100 ;
        RECT 39.800 111.100 40.200 113.000 ;
        RECT 41.400 111.100 41.800 113.000 ;
        RECT 44.000 111.100 44.400 113.900 ;
        RECT 45.400 112.800 45.800 113.200 ;
        RECT 46.300 113.100 46.600 114.900 ;
        RECT 47.800 114.800 50.600 114.900 ;
        RECT 47.000 113.800 47.400 114.600 ;
        RECT 45.500 112.400 45.900 112.800 ;
        RECT 46.200 111.100 46.600 113.100 ;
        RECT 50.200 111.100 50.600 114.800 ;
        RECT 52.600 115.100 53.000 119.900 ;
        RECT 54.500 119.200 54.900 119.900 ;
        RECT 54.500 118.800 55.400 119.200 ;
        RECT 53.400 115.800 53.800 116.600 ;
        RECT 54.500 116.300 54.900 118.800 ;
        RECT 54.500 115.900 55.400 116.300 ;
        RECT 54.200 115.100 54.600 115.600 ;
        RECT 52.600 114.800 54.600 115.100 ;
        RECT 51.800 113.400 52.200 114.200 ;
        RECT 51.000 112.400 51.400 113.200 ;
        RECT 52.600 113.100 53.000 114.800 ;
        RECT 55.000 114.200 55.300 115.900 ;
        RECT 56.600 115.600 57.000 119.900 ;
        RECT 58.700 119.200 59.100 119.900 ;
        RECT 58.700 118.800 59.400 119.200 ;
        RECT 58.700 116.200 59.100 118.800 ;
        RECT 58.700 115.900 59.400 116.200 ;
        RECT 59.800 115.900 60.200 119.900 ;
        RECT 60.600 116.200 61.000 119.900 ;
        RECT 62.200 116.200 62.600 119.900 ;
        RECT 60.600 115.900 62.600 116.200 ;
        RECT 56.600 115.400 58.600 115.600 ;
        RECT 56.600 115.300 58.700 115.400 ;
        RECT 58.300 115.000 58.700 115.300 ;
        RECT 59.100 115.200 59.400 115.900 ;
        RECT 59.900 115.200 60.200 115.900 ;
        RECT 61.800 115.200 62.200 115.400 ;
        RECT 57.600 114.200 58.000 114.600 ;
        RECT 54.200 113.800 54.600 114.200 ;
        RECT 55.000 113.800 55.400 114.200 ;
        RECT 57.400 114.100 57.900 114.200 ;
        RECT 55.800 113.800 57.900 114.100 ;
        RECT 54.200 113.100 54.500 113.800 ;
        RECT 52.600 112.800 54.500 113.100 ;
        RECT 53.100 111.100 53.500 112.800 ;
        RECT 55.000 112.100 55.300 113.800 ;
        RECT 55.800 113.200 56.100 113.800 ;
        RECT 58.400 113.500 58.700 115.000 ;
        RECT 59.000 114.800 59.400 115.200 ;
        RECT 59.800 114.900 61.000 115.200 ;
        RECT 61.800 115.100 62.600 115.200 ;
        RECT 63.000 115.100 63.400 119.900 ;
        RECT 64.600 115.900 65.000 119.900 ;
        RECT 65.400 116.200 65.800 119.900 ;
        RECT 67.000 116.200 67.400 119.900 ;
        RECT 68.600 117.900 69.000 119.900 ;
        RECT 68.700 117.800 69.000 117.900 ;
        RECT 70.200 117.900 70.600 119.900 ;
        RECT 70.200 117.800 70.500 117.900 ;
        RECT 68.700 117.500 70.500 117.800 ;
        RECT 69.400 116.400 69.800 117.200 ;
        RECT 70.200 116.200 70.500 117.500 ;
        RECT 72.300 117.200 72.700 119.900 ;
        RECT 74.200 117.900 74.600 119.900 ;
        RECT 74.300 117.800 74.600 117.900 ;
        RECT 75.800 117.900 76.200 119.900 ;
        RECT 75.800 117.800 76.100 117.900 ;
        RECT 74.300 117.500 76.100 117.800 ;
        RECT 71.800 116.800 72.700 117.200 ;
        RECT 73.000 116.800 73.400 117.200 ;
        RECT 72.300 116.200 72.700 116.800 ;
        RECT 73.100 116.200 73.400 116.800 ;
        RECT 74.300 116.200 74.600 117.500 ;
        RECT 75.000 116.400 75.400 117.200 ;
        RECT 65.400 115.900 67.400 116.200 ;
        RECT 64.700 115.200 65.000 115.900 ;
        RECT 67.800 115.400 68.200 116.200 ;
        RECT 70.200 115.800 70.600 116.200 ;
        RECT 72.300 115.900 72.800 116.200 ;
        RECT 73.100 115.900 73.800 116.200 ;
        RECT 66.600 115.200 67.000 115.400 ;
        RECT 61.800 114.900 63.400 115.100 ;
        RECT 59.800 114.800 60.200 114.900 ;
        RECT 57.500 113.200 58.700 113.500 ;
        RECT 55.800 112.400 56.200 113.200 ;
        RECT 56.600 112.400 57.000 113.200 ;
        RECT 57.500 112.100 57.800 113.200 ;
        RECT 59.100 113.100 59.400 114.800 ;
        RECT 59.800 114.100 60.200 114.200 ;
        RECT 60.700 114.100 61.000 114.900 ;
        RECT 62.200 114.800 63.400 114.900 ;
        RECT 64.600 114.900 65.800 115.200 ;
        RECT 66.600 114.900 67.400 115.200 ;
        RECT 64.600 114.800 65.000 114.900 ;
        RECT 59.800 113.800 61.000 114.100 ;
        RECT 61.400 113.800 61.800 114.600 ;
        RECT 55.000 111.100 55.400 112.100 ;
        RECT 57.400 111.100 57.800 112.100 ;
        RECT 59.000 111.100 59.400 113.100 ;
        RECT 59.800 112.800 60.200 113.200 ;
        RECT 60.700 113.100 61.000 113.800 ;
        RECT 59.900 112.400 60.300 112.800 ;
        RECT 60.600 111.100 61.000 113.100 ;
        RECT 63.000 111.100 63.400 114.800 ;
        RECT 63.800 113.400 64.200 114.200 ;
        RECT 64.600 112.800 65.000 113.200 ;
        RECT 65.500 113.100 65.800 114.900 ;
        RECT 67.000 114.800 67.400 114.900 ;
        RECT 68.600 114.800 69.400 115.200 ;
        RECT 70.200 115.100 70.500 115.800 ;
        RECT 71.000 115.100 71.400 115.200 ;
        RECT 70.200 114.800 71.400 115.100 ;
        RECT 66.200 113.800 66.600 114.600 ;
        RECT 70.200 114.200 70.500 114.800 ;
        RECT 71.800 114.400 72.200 115.200 ;
        RECT 72.500 114.200 72.800 115.900 ;
        RECT 73.400 115.800 73.800 115.900 ;
        RECT 74.200 115.800 74.600 116.200 ;
        RECT 74.300 114.200 74.600 115.800 ;
        RECT 76.600 115.400 77.000 116.200 ;
        RECT 75.400 114.800 76.200 115.200 ;
        RECT 69.700 114.100 70.500 114.200 ;
        RECT 69.600 113.900 70.500 114.100 ;
        RECT 71.000 114.100 71.400 114.200 ;
        RECT 64.700 112.400 65.100 112.800 ;
        RECT 65.400 111.100 65.800 113.100 ;
        RECT 69.600 111.100 70.000 113.900 ;
        RECT 71.000 113.800 71.800 114.100 ;
        RECT 72.500 113.800 73.800 114.200 ;
        RECT 74.300 114.100 75.100 114.200 ;
        RECT 78.200 114.100 78.600 119.900 ;
        RECT 80.300 116.200 80.700 119.900 ;
        RECT 83.000 118.200 83.400 119.900 ;
        RECT 82.900 117.900 83.400 118.200 ;
        RECT 82.900 117.600 83.200 117.900 ;
        RECT 84.600 117.600 85.000 119.900 ;
        RECT 86.200 118.500 86.600 119.900 ;
        RECT 87.000 118.500 87.400 119.900 ;
        RECT 82.200 117.300 83.200 117.600 ;
        RECT 81.000 116.800 81.400 117.200 ;
        RECT 81.100 116.200 81.400 116.800 ;
        RECT 80.300 115.900 80.800 116.200 ;
        RECT 81.100 115.900 81.800 116.200 ;
        RECT 80.500 115.200 80.800 115.900 ;
        RECT 81.400 115.800 81.800 115.900 ;
        RECT 79.000 115.100 79.400 115.200 ;
        RECT 79.800 115.100 80.200 115.200 ;
        RECT 79.000 114.800 80.200 115.100 ;
        RECT 79.800 114.400 80.200 114.800 ;
        RECT 80.500 114.800 81.000 115.200 ;
        RECT 80.500 114.200 80.800 114.800 ;
        RECT 82.200 114.500 82.600 117.300 ;
        RECT 83.500 117.200 85.600 117.600 ;
        RECT 87.800 117.500 88.200 119.900 ;
        RECT 89.400 117.500 89.800 119.900 ;
        RECT 83.500 117.000 83.800 117.200 ;
        RECT 83.000 116.600 83.800 117.000 ;
        RECT 85.300 116.900 88.200 117.200 ;
        RECT 84.300 116.600 85.000 116.900 ;
        RECT 84.300 116.500 87.400 116.600 ;
        RECT 84.700 116.300 87.400 116.500 ;
        RECT 87.000 116.200 87.400 116.300 ;
        RECT 87.900 116.500 88.200 116.900 ;
        RECT 88.500 116.800 89.800 117.200 ;
        RECT 91.000 116.800 91.400 119.900 ;
        RECT 91.800 118.500 92.200 119.900 ;
        RECT 92.600 118.500 93.000 119.900 ;
        RECT 93.400 118.500 93.800 119.900 ;
        RECT 92.600 117.200 94.700 117.600 ;
        RECT 95.000 117.200 95.400 119.900 ;
        RECT 96.600 117.600 97.000 119.900 ;
        RECT 96.600 117.300 97.900 117.600 ;
        RECT 95.000 116.800 96.300 117.200 ;
        RECT 91.800 116.500 92.200 116.600 ;
        RECT 87.900 116.200 92.200 116.500 ;
        RECT 93.400 116.500 93.800 116.600 ;
        RECT 97.600 116.500 97.900 117.300 ;
        RECT 93.400 116.200 97.900 116.500 ;
        RECT 97.600 115.300 97.900 116.200 ;
        RECT 98.200 116.000 98.600 119.900 ;
        RECT 101.700 117.200 102.100 119.900 ;
        RECT 101.700 116.800 102.600 117.200 ;
        RECT 101.700 116.300 102.100 116.800 ;
        RECT 98.200 115.600 98.700 116.000 ;
        RECT 101.700 115.900 102.600 116.300 ;
        RECT 82.900 115.000 94.600 115.300 ;
        RECT 97.600 115.000 98.000 115.300 ;
        RECT 82.900 114.900 83.300 115.000 ;
        RECT 84.600 114.800 85.000 115.000 ;
        RECT 85.400 114.800 85.800 115.000 ;
        RECT 94.200 114.700 94.600 115.000 ;
        RECT 79.000 114.100 79.400 114.200 ;
        RECT 74.300 113.900 75.200 114.100 ;
        RECT 71.400 113.600 71.800 113.800 ;
        RECT 71.100 113.100 72.900 113.300 ;
        RECT 73.400 113.100 73.700 113.800 ;
        RECT 71.000 113.000 73.000 113.100 ;
        RECT 71.000 111.100 71.400 113.000 ;
        RECT 72.600 111.100 73.000 113.000 ;
        RECT 73.400 111.100 73.800 113.100 ;
        RECT 74.800 111.100 75.200 113.900 ;
        RECT 78.200 113.800 79.800 114.100 ;
        RECT 80.500 113.800 81.800 114.200 ;
        RECT 82.200 114.100 86.600 114.500 ;
        RECT 86.900 114.300 87.900 114.700 ;
        RECT 89.800 114.300 91.400 114.700 ;
        RECT 77.400 112.400 77.800 113.200 ;
        RECT 78.200 111.100 78.600 113.800 ;
        RECT 79.400 113.600 79.800 113.800 ;
        RECT 79.100 113.100 80.900 113.300 ;
        RECT 81.400 113.100 81.700 113.800 ;
        RECT 79.000 113.000 81.000 113.100 ;
        RECT 79.000 111.100 79.400 113.000 ;
        RECT 80.600 111.100 81.000 113.000 ;
        RECT 81.400 111.100 81.800 113.100 ;
        RECT 82.200 111.100 82.600 114.100 ;
        RECT 83.400 113.400 84.900 113.800 ;
        RECT 84.500 113.100 84.900 113.400 ;
        RECT 87.500 113.100 87.900 114.300 ;
        RECT 88.600 113.400 89.000 114.200 ;
        RECT 91.200 113.900 91.600 114.000 ;
        RECT 89.400 113.600 91.600 113.900 ;
        RECT 89.400 113.500 89.800 113.600 ;
        RECT 92.600 113.200 93.000 114.600 ;
        RECT 95.500 114.300 97.400 114.700 ;
        RECT 95.500 113.700 95.900 114.300 ;
        RECT 97.700 114.000 98.000 115.000 ;
        RECT 89.400 113.100 89.800 113.200 ;
        RECT 84.500 112.700 85.800 113.100 ;
        RECT 87.500 112.800 89.800 113.100 ;
        RECT 92.500 112.800 93.000 113.200 ;
        RECT 95.000 113.400 95.900 113.700 ;
        RECT 97.400 113.700 98.000 114.000 ;
        RECT 95.000 113.100 95.400 113.400 ;
        RECT 85.400 111.100 85.800 112.700 ;
        RECT 94.200 112.700 95.400 113.100 ;
        RECT 86.200 111.100 86.600 112.500 ;
        RECT 87.000 111.100 87.400 112.500 ;
        RECT 87.800 111.100 88.200 112.500 ;
        RECT 89.400 111.100 89.800 112.500 ;
        RECT 91.000 111.100 91.400 112.500 ;
        RECT 91.800 111.100 92.200 112.500 ;
        RECT 92.600 111.100 93.000 112.500 ;
        RECT 93.400 111.100 93.800 112.500 ;
        RECT 94.200 111.100 94.600 112.700 ;
        RECT 97.400 111.100 97.800 113.700 ;
        RECT 98.300 113.400 98.700 115.600 ;
        RECT 99.800 115.100 100.200 115.200 ;
        RECT 101.400 115.100 101.800 115.600 ;
        RECT 99.800 114.800 101.800 115.100 ;
        RECT 98.200 113.000 98.700 113.400 ;
        RECT 102.200 114.200 102.500 115.900 ;
        RECT 102.200 113.800 102.600 114.200 ;
        RECT 104.600 114.100 105.000 119.900 ;
        RECT 105.400 119.600 107.400 119.900 ;
        RECT 105.400 115.900 105.800 119.600 ;
        RECT 106.200 115.900 106.600 119.300 ;
        RECT 107.000 116.200 107.400 119.600 ;
        RECT 108.600 116.200 109.000 119.900 ;
        RECT 109.400 117.900 109.800 119.900 ;
        RECT 109.500 117.800 109.800 117.900 ;
        RECT 111.000 117.900 111.400 119.900 ;
        RECT 111.000 117.800 111.300 117.900 ;
        RECT 109.500 117.500 111.300 117.800 ;
        RECT 109.500 116.200 109.800 117.500 ;
        RECT 110.200 116.400 110.600 117.200 ;
        RECT 111.000 117.100 111.400 117.200 ;
        RECT 112.600 117.100 113.000 119.900 ;
        RECT 111.000 116.800 113.000 117.100 ;
        RECT 107.000 115.900 109.000 116.200 ;
        RECT 106.300 115.600 106.600 115.900 ;
        RECT 109.400 115.800 109.800 116.200 ;
        RECT 105.400 114.800 105.800 115.600 ;
        RECT 106.300 115.300 107.300 115.600 ;
        RECT 107.000 115.200 107.300 115.300 ;
        RECT 108.200 115.200 108.600 115.400 ;
        RECT 107.000 114.800 107.400 115.200 ;
        RECT 108.200 114.900 109.000 115.200 ;
        RECT 108.600 114.800 109.000 114.900 ;
        RECT 106.300 114.400 106.700 114.800 ;
        RECT 106.300 114.200 106.600 114.400 ;
        RECT 105.400 114.100 105.800 114.200 ;
        RECT 104.600 113.800 105.800 114.100 ;
        RECT 106.200 113.800 106.600 114.200 ;
        RECT 98.200 111.100 98.600 113.000 ;
        RECT 102.200 112.100 102.500 113.800 ;
        RECT 103.000 112.400 103.400 113.200 ;
        RECT 102.200 111.100 102.600 112.100 ;
        RECT 104.600 111.100 105.000 113.800 ;
        RECT 107.000 113.100 107.300 114.800 ;
        RECT 107.800 113.800 108.200 114.600 ;
        RECT 109.500 114.200 109.800 115.800 ;
        RECT 111.800 115.400 112.200 116.200 ;
        RECT 110.600 114.800 111.400 115.200 ;
        RECT 109.500 114.100 110.300 114.200 ;
        RECT 109.500 113.900 110.400 114.100 ;
        RECT 106.700 111.100 107.500 113.100 ;
        RECT 110.000 112.100 110.400 113.900 ;
        RECT 111.000 112.100 111.400 112.200 ;
        RECT 110.000 111.800 111.400 112.100 ;
        RECT 110.000 111.100 110.400 111.800 ;
        RECT 112.600 111.100 113.000 116.800 ;
        RECT 114.200 116.200 114.600 119.900 ;
        RECT 115.800 119.600 117.800 119.900 ;
        RECT 115.800 116.200 116.200 119.600 ;
        RECT 114.200 115.900 116.200 116.200 ;
        RECT 116.600 115.900 117.000 119.300 ;
        RECT 117.400 115.900 117.800 119.600 ;
        RECT 118.200 116.200 118.600 119.900 ;
        RECT 119.800 119.600 121.800 119.900 ;
        RECT 119.800 116.200 120.200 119.600 ;
        RECT 118.200 115.900 120.200 116.200 ;
        RECT 116.600 115.600 116.900 115.900 ;
        RECT 120.600 115.800 121.000 119.300 ;
        RECT 121.400 115.900 121.800 119.600 ;
        RECT 123.000 118.200 123.400 119.900 ;
        RECT 122.900 117.900 123.400 118.200 ;
        RECT 122.900 117.600 123.200 117.900 ;
        RECT 124.600 117.600 125.000 119.900 ;
        RECT 126.200 118.500 126.600 119.900 ;
        RECT 127.000 118.500 127.400 119.900 ;
        RECT 122.200 117.300 123.200 117.600 ;
        RECT 120.600 115.600 120.900 115.800 ;
        RECT 114.600 115.200 115.000 115.400 ;
        RECT 115.900 115.300 116.900 115.600 ;
        RECT 115.900 115.200 116.200 115.300 ;
        RECT 114.200 114.900 115.000 115.200 ;
        RECT 114.200 114.800 114.600 114.900 ;
        RECT 115.800 114.800 116.200 115.200 ;
        RECT 117.400 114.800 117.800 115.600 ;
        RECT 118.600 115.200 119.000 115.400 ;
        RECT 119.900 115.300 120.900 115.600 ;
        RECT 119.900 115.200 120.200 115.300 ;
        RECT 118.200 114.900 119.000 115.200 ;
        RECT 118.200 114.800 118.600 114.900 ;
        RECT 119.800 114.800 120.200 115.200 ;
        RECT 121.400 114.800 121.800 115.600 ;
        RECT 115.000 113.800 115.400 114.600 ;
        RECT 113.400 112.400 113.800 113.200 ;
        RECT 115.900 113.100 116.200 114.800 ;
        RECT 116.500 114.400 116.900 114.800 ;
        RECT 116.600 114.200 116.900 114.400 ;
        RECT 117.400 114.200 117.700 114.800 ;
        RECT 116.600 113.800 117.000 114.200 ;
        RECT 117.400 113.800 117.800 114.200 ;
        RECT 119.000 113.800 119.400 114.600 ;
        RECT 119.900 113.100 120.200 114.800 ;
        RECT 120.500 114.400 120.900 114.800 ;
        RECT 120.600 114.200 120.900 114.400 ;
        RECT 122.200 114.500 122.600 117.300 ;
        RECT 123.500 117.200 125.600 117.600 ;
        RECT 127.800 117.500 128.200 119.900 ;
        RECT 129.400 117.500 129.800 119.900 ;
        RECT 123.500 117.000 123.800 117.200 ;
        RECT 123.000 116.600 123.800 117.000 ;
        RECT 125.300 116.900 128.200 117.200 ;
        RECT 124.300 116.600 125.000 116.900 ;
        RECT 124.300 116.500 127.400 116.600 ;
        RECT 124.700 116.300 127.400 116.500 ;
        RECT 127.000 116.200 127.400 116.300 ;
        RECT 127.900 116.500 128.200 116.900 ;
        RECT 128.500 116.800 129.800 117.200 ;
        RECT 131.000 116.800 131.400 119.900 ;
        RECT 131.800 118.500 132.200 119.900 ;
        RECT 132.600 118.500 133.000 119.900 ;
        RECT 133.400 118.500 133.800 119.900 ;
        RECT 132.600 117.200 134.700 117.600 ;
        RECT 135.000 117.200 135.400 119.900 ;
        RECT 136.600 117.600 137.000 119.900 ;
        RECT 136.600 117.300 137.900 117.600 ;
        RECT 135.000 116.800 136.300 117.200 ;
        RECT 131.800 116.500 132.200 116.600 ;
        RECT 127.900 116.200 132.200 116.500 ;
        RECT 133.400 116.500 133.800 116.600 ;
        RECT 137.600 116.500 137.900 117.300 ;
        RECT 133.400 116.200 137.900 116.500 ;
        RECT 137.600 115.300 137.900 116.200 ;
        RECT 138.200 116.000 138.600 119.900 ;
        RECT 138.200 115.600 138.700 116.000 ;
        RECT 122.900 115.000 134.600 115.300 ;
        RECT 137.600 115.000 138.000 115.300 ;
        RECT 122.900 114.900 123.300 115.000 ;
        RECT 124.600 114.800 125.000 115.000 ;
        RECT 125.400 114.800 125.800 115.000 ;
        RECT 134.200 114.700 134.600 115.000 ;
        RECT 120.600 113.800 121.000 114.200 ;
        RECT 122.200 114.100 126.600 114.500 ;
        RECT 126.900 114.300 127.900 114.700 ;
        RECT 129.800 114.300 131.400 114.700 ;
        RECT 115.700 111.100 116.500 113.100 ;
        RECT 119.700 111.100 120.500 113.100 ;
        RECT 122.200 111.100 122.600 114.100 ;
        RECT 123.400 113.400 124.900 113.800 ;
        RECT 124.500 113.100 124.900 113.400 ;
        RECT 127.500 113.100 127.900 114.300 ;
        RECT 128.600 113.400 129.000 114.200 ;
        RECT 131.200 113.900 131.600 114.000 ;
        RECT 129.400 113.600 131.600 113.900 ;
        RECT 129.400 113.500 129.800 113.600 ;
        RECT 132.600 113.200 133.000 114.600 ;
        RECT 135.500 114.300 137.400 114.700 ;
        RECT 135.500 113.700 135.900 114.300 ;
        RECT 137.700 114.000 138.000 115.000 ;
        RECT 129.400 113.100 129.800 113.200 ;
        RECT 124.500 112.700 125.800 113.100 ;
        RECT 127.500 112.800 129.800 113.100 ;
        RECT 132.500 112.800 133.000 113.200 ;
        RECT 135.000 113.400 135.900 113.700 ;
        RECT 137.400 113.700 138.000 114.000 ;
        RECT 138.300 114.100 138.700 115.600 ;
        RECT 139.000 114.100 139.400 114.200 ;
        RECT 138.300 113.800 139.400 114.100 ;
        RECT 135.000 113.100 135.400 113.400 ;
        RECT 125.400 111.100 125.800 112.700 ;
        RECT 134.200 112.700 135.400 113.100 ;
        RECT 126.200 111.100 126.600 112.500 ;
        RECT 127.000 111.100 127.400 112.500 ;
        RECT 127.800 111.100 128.200 112.500 ;
        RECT 129.400 111.100 129.800 112.500 ;
        RECT 131.000 111.100 131.400 112.500 ;
        RECT 131.800 111.100 132.200 112.500 ;
        RECT 132.600 111.100 133.000 112.500 ;
        RECT 133.400 111.100 133.800 112.500 ;
        RECT 134.200 111.100 134.600 112.700 ;
        RECT 137.400 111.100 137.800 113.700 ;
        RECT 138.300 113.400 138.700 113.800 ;
        RECT 138.200 113.000 138.700 113.400 ;
        RECT 138.200 111.100 138.600 113.000 ;
        RECT 139.800 111.100 140.200 119.900 ;
        RECT 141.400 116.200 141.800 119.900 ;
        RECT 143.800 116.200 144.200 119.900 ;
        RECT 146.200 116.200 146.600 119.900 ;
        RECT 141.400 115.900 142.500 116.200 ;
        RECT 143.800 115.900 144.900 116.200 ;
        RECT 146.200 115.900 147.300 116.200 ;
        RECT 142.200 115.600 142.500 115.900 ;
        RECT 144.600 115.600 144.900 115.900 ;
        RECT 147.000 115.600 147.300 115.900 ;
        RECT 142.200 115.200 142.800 115.600 ;
        RECT 144.600 115.200 145.200 115.600 ;
        RECT 147.000 115.200 147.600 115.600 ;
        RECT 140.600 115.100 141.000 115.200 ;
        RECT 141.400 115.100 141.800 115.200 ;
        RECT 140.600 114.800 141.800 115.100 ;
        RECT 141.400 114.400 141.800 114.800 ;
        RECT 142.200 113.700 142.500 115.200 ;
        RECT 143.800 114.400 144.200 115.200 ;
        RECT 144.600 113.700 144.900 115.200 ;
        RECT 146.200 114.400 146.600 115.200 ;
        RECT 147.000 113.700 147.300 115.200 ;
        RECT 141.400 113.400 142.500 113.700 ;
        RECT 143.800 113.400 144.900 113.700 ;
        RECT 146.200 113.400 147.300 113.700 ;
        RECT 140.600 112.400 141.000 113.200 ;
        RECT 141.400 111.100 141.800 113.400 ;
        RECT 143.800 111.100 144.200 113.400 ;
        RECT 146.200 111.100 146.600 113.400 ;
        RECT 0.600 107.900 1.000 109.900 ;
        RECT 1.400 108.000 1.800 109.900 ;
        RECT 3.000 108.000 3.400 109.900 ;
        RECT 3.900 108.200 4.300 108.600 ;
        RECT 1.400 107.900 3.400 108.000 ;
        RECT 0.700 107.200 1.000 107.900 ;
        RECT 1.500 107.700 3.300 107.900 ;
        RECT 3.800 107.800 4.200 108.200 ;
        RECT 4.600 107.900 5.000 109.900 ;
        RECT 2.600 107.200 3.000 107.400 ;
        RECT 0.600 106.800 1.900 107.200 ;
        RECT 2.600 107.100 3.400 107.200 ;
        RECT 4.700 107.100 5.000 107.900 ;
        RECT 2.600 106.900 5.000 107.100 ;
        RECT 3.000 106.800 5.000 106.900 ;
        RECT 0.600 105.100 1.000 105.200 ;
        RECT 1.600 105.100 1.900 106.800 ;
        RECT 2.200 106.100 2.600 106.600 ;
        RECT 3.000 106.100 3.400 106.200 ;
        RECT 2.200 105.800 3.400 106.100 ;
        RECT 3.800 106.100 4.200 106.200 ;
        RECT 4.700 106.100 5.000 106.800 ;
        RECT 5.400 106.400 5.800 107.200 ;
        RECT 7.600 107.100 8.000 109.900 ;
        RECT 7.100 106.900 8.000 107.100 ;
        RECT 12.000 107.100 12.400 109.900 ;
        RECT 14.700 108.200 15.100 109.900 ;
        RECT 14.200 107.900 15.100 108.200 ;
        RECT 12.000 106.900 12.900 107.100 ;
        RECT 7.100 106.800 7.900 106.900 ;
        RECT 12.100 106.800 12.900 106.900 ;
        RECT 13.400 106.800 13.800 107.600 ;
        RECT 6.200 106.100 6.600 106.200 ;
        RECT 3.800 105.800 5.000 106.100 ;
        RECT 5.800 105.800 6.600 106.100 ;
        RECT 3.900 105.100 4.200 105.800 ;
        RECT 5.800 105.600 6.200 105.800 ;
        RECT 7.100 105.200 7.400 106.800 ;
        RECT 8.200 105.800 9.000 106.200 ;
        RECT 11.000 105.800 11.800 106.200 ;
        RECT 0.600 104.800 1.300 105.100 ;
        RECT 1.600 104.800 2.100 105.100 ;
        RECT 1.000 104.200 1.300 104.800 ;
        RECT 1.700 104.200 2.100 104.800 ;
        RECT 1.000 103.800 1.400 104.200 ;
        RECT 1.700 103.800 2.600 104.200 ;
        RECT 1.700 101.100 2.100 103.800 ;
        RECT 3.800 101.100 4.200 105.100 ;
        RECT 4.600 104.800 6.600 105.100 ;
        RECT 7.000 104.800 7.400 105.200 ;
        RECT 9.400 105.100 9.800 105.600 ;
        RECT 10.200 105.100 10.600 105.600 ;
        RECT 9.400 104.800 10.600 105.100 ;
        RECT 12.600 105.200 12.900 106.800 ;
        RECT 12.600 104.800 13.000 105.200 ;
        RECT 4.600 101.100 5.000 104.800 ;
        RECT 6.200 101.100 6.600 104.800 ;
        RECT 7.100 103.500 7.400 104.800 ;
        RECT 7.800 104.100 8.200 104.600 ;
        RECT 11.800 104.100 12.200 104.600 ;
        RECT 7.800 103.800 12.200 104.100 ;
        RECT 12.600 103.500 12.900 104.800 ;
        RECT 7.100 103.200 8.900 103.500 ;
        RECT 7.100 103.100 7.400 103.200 ;
        RECT 7.000 101.100 7.400 103.100 ;
        RECT 8.600 103.100 8.900 103.200 ;
        RECT 11.100 103.200 12.900 103.500 ;
        RECT 11.100 103.100 11.400 103.200 ;
        RECT 8.600 101.100 9.000 103.100 ;
        RECT 11.000 101.100 11.400 103.100 ;
        RECT 12.600 103.100 12.900 103.200 ;
        RECT 12.600 101.100 13.000 103.100 ;
        RECT 14.200 101.100 14.600 107.900 ;
        RECT 15.800 106.800 16.200 107.600 ;
        RECT 16.600 107.100 17.000 109.900 ;
        RECT 18.700 108.200 19.100 109.900 ;
        RECT 18.200 107.900 19.100 108.200 ;
        RECT 17.400 107.100 17.800 107.600 ;
        RECT 16.600 106.800 17.800 107.100 ;
        RECT 15.000 104.400 15.400 105.200 ;
        RECT 16.600 101.100 17.000 106.800 ;
        RECT 18.200 101.100 18.600 107.900 ;
        RECT 20.400 107.100 20.800 109.900 ;
        RECT 23.600 107.100 24.000 109.900 ;
        RECT 26.300 108.200 26.700 108.600 ;
        RECT 24.600 107.800 25.000 108.200 ;
        RECT 26.200 107.800 26.600 108.200 ;
        RECT 27.000 107.900 27.400 109.900 ;
        RECT 30.200 109.100 30.600 109.200 ;
        RECT 31.200 109.100 31.600 109.900 ;
        RECT 30.200 108.800 31.600 109.100 ;
        RECT 24.600 107.100 24.900 107.800 ;
        RECT 19.900 106.900 20.800 107.100 ;
        RECT 19.900 106.800 20.700 106.900 ;
        RECT 23.100 106.800 24.900 107.100 ;
        RECT 19.900 105.200 20.200 106.800 ;
        RECT 21.000 105.800 21.800 106.200 ;
        RECT 19.000 104.400 19.400 105.200 ;
        RECT 19.800 104.800 20.200 105.200 ;
        RECT 22.200 104.800 22.600 105.600 ;
        RECT 23.100 105.200 23.400 106.800 ;
        RECT 24.200 105.800 25.000 106.200 ;
        RECT 23.000 104.800 23.400 105.200 ;
        RECT 25.400 104.800 25.800 106.200 ;
        RECT 26.200 106.100 26.600 106.200 ;
        RECT 27.100 106.100 27.400 107.900 ;
        RECT 27.800 106.400 28.200 107.200 ;
        RECT 31.200 107.100 31.600 108.800 ;
        RECT 34.400 107.100 34.800 109.900 ;
        RECT 35.900 108.200 36.300 108.600 ;
        RECT 35.800 107.800 36.200 108.200 ;
        RECT 36.600 107.900 37.000 109.900 ;
        RECT 39.100 108.200 39.500 108.600 ;
        RECT 31.200 106.900 32.100 107.100 ;
        RECT 34.400 106.900 35.300 107.100 ;
        RECT 31.300 106.800 32.100 106.900 ;
        RECT 34.500 106.800 35.300 106.900 ;
        RECT 28.600 106.100 29.000 106.200 ;
        RECT 26.200 105.800 27.400 106.100 ;
        RECT 28.200 105.800 29.800 106.100 ;
        RECT 30.200 105.800 31.000 106.200 ;
        RECT 26.300 105.100 26.600 105.800 ;
        RECT 28.200 105.600 28.600 105.800 ;
        RECT 19.900 103.500 20.200 104.800 ;
        RECT 20.600 103.800 21.000 104.600 ;
        RECT 23.100 103.500 23.400 104.800 ;
        RECT 23.800 103.800 24.200 104.600 ;
        RECT 19.900 103.200 21.700 103.500 ;
        RECT 23.100 103.200 24.900 103.500 ;
        RECT 19.900 103.100 20.200 103.200 ;
        RECT 19.800 101.100 20.200 103.100 ;
        RECT 21.400 101.100 21.800 103.200 ;
        RECT 23.100 103.100 23.400 103.200 ;
        RECT 23.000 101.100 23.400 103.100 ;
        RECT 24.600 103.100 24.900 103.200 ;
        RECT 24.600 101.100 25.000 103.100 ;
        RECT 26.200 101.100 26.600 105.100 ;
        RECT 27.000 104.800 29.000 105.100 ;
        RECT 29.400 104.800 29.800 105.800 ;
        RECT 31.800 105.200 32.100 106.800 ;
        RECT 33.400 105.800 34.200 106.200 ;
        RECT 31.800 104.800 32.200 105.200 ;
        RECT 32.600 104.800 33.000 105.600 ;
        RECT 35.000 105.200 35.300 106.800 ;
        RECT 35.800 106.100 36.200 106.200 ;
        RECT 36.700 106.100 37.000 107.900 ;
        RECT 39.000 107.800 39.400 108.200 ;
        RECT 39.800 107.900 40.200 109.900 ;
        RECT 43.000 109.100 43.400 109.200 ;
        RECT 44.000 109.100 44.400 109.900 ;
        RECT 43.000 108.800 44.400 109.100 ;
        RECT 37.400 106.400 37.800 107.200 ;
        RECT 38.200 106.100 38.600 106.200 ;
        RECT 35.800 105.800 37.000 106.100 ;
        RECT 37.800 105.800 38.600 106.100 ;
        RECT 39.000 106.100 39.400 106.200 ;
        RECT 39.900 106.100 40.200 107.900 ;
        RECT 40.600 106.400 41.000 107.200 ;
        RECT 44.000 107.100 44.400 108.800 ;
        RECT 47.200 107.100 47.600 109.900 ;
        RECT 52.000 109.200 52.400 109.900 ;
        RECT 51.800 108.800 52.400 109.200 ;
        RECT 52.000 107.100 52.400 108.800 ;
        RECT 53.400 107.900 53.800 109.900 ;
        RECT 54.200 108.000 54.600 109.900 ;
        RECT 55.800 108.000 56.200 109.900 ;
        RECT 54.200 107.900 56.200 108.000 ;
        RECT 56.600 107.900 57.000 109.900 ;
        RECT 57.400 108.000 57.800 109.900 ;
        RECT 59.000 108.000 59.400 109.900 ;
        RECT 57.400 107.900 59.400 108.000 ;
        RECT 61.400 107.900 61.800 109.900 ;
        RECT 62.100 108.200 62.500 108.600 ;
        RECT 53.500 107.200 53.800 107.900 ;
        RECT 54.300 107.700 56.100 107.900 ;
        RECT 55.400 107.200 55.800 107.400 ;
        RECT 56.700 107.200 57.000 107.900 ;
        RECT 57.500 107.700 59.300 107.900 ;
        RECT 58.600 107.200 59.000 107.400 ;
        RECT 44.000 106.900 44.900 107.100 ;
        RECT 47.200 106.900 48.100 107.100 ;
        RECT 52.000 106.900 52.900 107.100 ;
        RECT 44.100 106.800 44.900 106.900 ;
        RECT 47.300 106.800 48.100 106.900 ;
        RECT 52.100 106.800 52.900 106.900 ;
        RECT 53.400 106.800 54.700 107.200 ;
        RECT 55.400 106.900 56.200 107.200 ;
        RECT 55.800 106.800 56.200 106.900 ;
        RECT 56.600 106.800 57.900 107.200 ;
        RECT 58.600 106.900 59.400 107.200 ;
        RECT 59.000 106.800 59.400 106.900 ;
        RECT 41.400 106.100 41.800 106.200 ;
        RECT 39.000 105.800 40.200 106.100 ;
        RECT 41.000 105.800 42.600 106.100 ;
        RECT 43.000 105.800 43.800 106.200 ;
        RECT 35.000 104.800 35.400 105.200 ;
        RECT 35.900 105.100 36.200 105.800 ;
        RECT 37.800 105.600 38.200 105.800 ;
        RECT 39.100 105.100 39.400 105.800 ;
        RECT 41.000 105.600 41.400 105.800 ;
        RECT 27.000 101.100 27.400 104.800 ;
        RECT 28.600 101.100 29.000 104.800 ;
        RECT 31.000 103.800 31.400 104.600 ;
        RECT 31.800 103.500 32.100 104.800 ;
        RECT 34.200 103.800 34.600 104.600 ;
        RECT 35.000 103.500 35.300 104.800 ;
        RECT 30.300 103.200 32.100 103.500 ;
        RECT 30.300 103.100 30.600 103.200 ;
        RECT 30.200 101.100 30.600 103.100 ;
        RECT 31.800 103.100 32.100 103.200 ;
        RECT 33.500 103.200 35.300 103.500 ;
        RECT 33.500 103.100 33.800 103.200 ;
        RECT 31.800 101.100 32.200 103.100 ;
        RECT 33.400 101.100 33.800 103.100 ;
        RECT 35.000 103.100 35.300 103.200 ;
        RECT 35.000 101.100 35.400 103.100 ;
        RECT 35.800 101.100 36.200 105.100 ;
        RECT 36.600 104.800 38.600 105.100 ;
        RECT 36.600 101.100 37.000 104.800 ;
        RECT 38.200 101.100 38.600 104.800 ;
        RECT 39.000 101.100 39.400 105.100 ;
        RECT 39.800 104.800 41.800 105.100 ;
        RECT 42.200 104.800 42.600 105.800 ;
        RECT 44.600 105.200 44.900 106.800 ;
        RECT 46.200 105.800 47.000 106.200 ;
        RECT 47.800 106.100 48.100 106.800 ;
        RECT 48.600 106.100 49.000 106.200 ;
        RECT 47.800 105.800 49.000 106.100 ;
        RECT 51.000 105.800 51.800 106.200 ;
        RECT 44.600 104.800 45.000 105.200 ;
        RECT 45.400 104.800 45.800 105.600 ;
        RECT 47.800 105.200 48.100 105.800 ;
        RECT 47.800 104.800 48.200 105.200 ;
        RECT 50.200 104.800 50.600 105.600 ;
        RECT 52.600 105.200 52.900 106.800 ;
        RECT 52.600 104.800 53.000 105.200 ;
        RECT 53.400 105.100 53.800 105.200 ;
        RECT 54.400 105.100 54.700 106.800 ;
        RECT 55.000 106.100 55.400 106.600 ;
        RECT 57.600 106.200 57.900 106.800 ;
        RECT 55.000 105.800 56.900 106.100 ;
        RECT 57.400 105.800 57.900 106.200 ;
        RECT 58.200 106.100 58.600 106.600 ;
        RECT 60.600 106.400 61.000 107.200 ;
        RECT 59.000 106.100 59.400 106.200 ;
        RECT 58.200 105.800 59.400 106.100 ;
        RECT 59.800 106.100 60.200 106.200 ;
        RECT 61.400 106.100 61.700 107.900 ;
        RECT 62.200 107.800 62.600 108.200 ;
        RECT 63.000 108.000 63.400 109.900 ;
        RECT 64.600 108.000 65.000 109.900 ;
        RECT 63.000 107.900 65.000 108.000 ;
        RECT 65.400 107.900 65.800 109.900 ;
        RECT 66.200 107.900 66.600 109.900 ;
        RECT 67.000 108.000 67.400 109.900 ;
        RECT 68.600 108.000 69.000 109.900 ;
        RECT 67.000 107.900 69.000 108.000 ;
        RECT 63.100 107.700 64.900 107.900 ;
        RECT 63.400 107.200 63.800 107.400 ;
        RECT 65.400 107.200 65.700 107.900 ;
        RECT 66.300 107.200 66.600 107.900 ;
        RECT 67.100 107.700 68.900 107.900 ;
        RECT 68.200 107.200 68.600 107.400 ;
        RECT 63.000 106.900 63.800 107.200 ;
        RECT 63.000 106.800 63.400 106.900 ;
        RECT 64.500 106.800 65.800 107.200 ;
        RECT 66.200 106.800 67.500 107.200 ;
        RECT 68.200 106.900 69.000 107.200 ;
        RECT 70.000 107.100 70.400 109.900 ;
        RECT 72.700 108.200 73.100 108.600 ;
        RECT 72.600 107.800 73.000 108.200 ;
        RECT 73.400 107.900 73.800 109.900 ;
        RECT 77.100 108.200 77.500 109.900 ;
        RECT 68.600 106.800 69.000 106.900 ;
        RECT 69.500 106.900 70.400 107.100 ;
        RECT 72.600 107.100 73.000 107.200 ;
        RECT 73.500 107.100 73.800 107.900 ;
        RECT 76.600 107.900 77.500 108.200 ;
        RECT 69.500 106.800 70.300 106.900 ;
        RECT 72.600 106.800 73.800 107.100 ;
        RECT 62.200 106.100 62.600 106.200 ;
        RECT 59.800 105.800 60.600 106.100 ;
        RECT 61.400 105.800 62.600 106.100 ;
        RECT 63.800 105.800 64.200 106.600 ;
        RECT 56.600 105.200 56.900 105.800 ;
        RECT 56.600 105.100 57.000 105.200 ;
        RECT 57.600 105.100 57.900 105.800 ;
        RECT 60.200 105.600 60.600 105.800 ;
        RECT 62.200 105.100 62.500 105.800 ;
        RECT 64.500 105.100 64.800 106.800 ;
        RECT 65.400 105.100 65.800 105.200 ;
        RECT 53.400 104.800 54.100 105.100 ;
        RECT 54.400 104.800 54.900 105.100 ;
        RECT 56.600 104.800 57.300 105.100 ;
        RECT 57.600 104.800 58.100 105.100 ;
        RECT 39.800 101.100 40.200 104.800 ;
        RECT 41.400 101.100 41.800 104.800 ;
        RECT 43.800 103.800 44.200 104.600 ;
        RECT 44.600 103.500 44.900 104.800 ;
        RECT 47.000 103.800 47.400 104.600 ;
        RECT 47.800 103.500 48.100 104.800 ;
        RECT 51.800 103.800 52.200 104.600 ;
        RECT 52.600 103.500 52.900 104.800 ;
        RECT 53.800 104.200 54.100 104.800 ;
        RECT 54.500 104.200 54.900 104.800 ;
        RECT 57.000 104.200 57.300 104.800 ;
        RECT 53.800 103.800 54.200 104.200 ;
        RECT 54.500 103.800 55.400 104.200 ;
        RECT 57.000 103.800 57.400 104.200 ;
        RECT 43.100 103.200 44.900 103.500 ;
        RECT 43.100 103.100 43.400 103.200 ;
        RECT 43.000 101.100 43.400 103.100 ;
        RECT 44.600 103.100 44.900 103.200 ;
        RECT 46.300 103.200 48.100 103.500 ;
        RECT 46.300 103.100 46.600 103.200 ;
        RECT 44.600 101.100 45.000 103.100 ;
        RECT 46.200 101.100 46.600 103.100 ;
        RECT 47.800 103.100 48.100 103.200 ;
        RECT 51.100 103.200 52.900 103.500 ;
        RECT 51.100 103.100 51.400 103.200 ;
        RECT 47.800 101.100 48.200 103.100 ;
        RECT 51.000 101.100 51.400 103.100 ;
        RECT 52.600 103.100 52.900 103.200 ;
        RECT 52.600 101.100 53.000 103.100 ;
        RECT 54.500 101.100 54.900 103.800 ;
        RECT 57.700 101.100 58.100 104.800 ;
        RECT 59.800 104.800 61.800 105.100 ;
        RECT 59.800 101.100 60.200 104.800 ;
        RECT 61.400 101.100 61.800 104.800 ;
        RECT 62.200 101.100 62.600 105.100 ;
        RECT 64.300 104.800 64.800 105.100 ;
        RECT 65.100 104.800 65.800 105.100 ;
        RECT 66.200 105.100 66.600 105.200 ;
        RECT 67.200 105.100 67.500 106.800 ;
        RECT 67.800 105.800 68.200 106.600 ;
        RECT 69.500 105.200 69.800 106.800 ;
        RECT 70.600 105.800 71.400 106.200 ;
        RECT 72.600 106.100 73.000 106.200 ;
        RECT 73.500 106.100 73.800 106.800 ;
        RECT 74.200 106.400 74.600 107.200 ;
        RECT 75.800 106.800 76.200 107.600 ;
        RECT 75.000 106.100 75.400 106.200 ;
        RECT 76.600 106.100 77.000 107.900 ;
        RECT 72.600 105.800 73.800 106.100 ;
        RECT 74.600 105.800 75.400 106.100 ;
        RECT 75.800 105.800 77.000 106.100 ;
        RECT 66.200 104.800 66.900 105.100 ;
        RECT 67.200 104.800 67.700 105.100 ;
        RECT 69.400 104.800 69.800 105.200 ;
        RECT 71.800 104.800 72.200 105.600 ;
        RECT 72.700 105.100 73.000 105.800 ;
        RECT 74.600 105.600 75.000 105.800 ;
        RECT 75.800 105.200 76.100 105.800 ;
        RECT 64.300 101.100 64.700 104.800 ;
        RECT 65.100 104.200 65.400 104.800 ;
        RECT 65.000 103.800 65.400 104.200 ;
        RECT 66.600 104.200 66.900 104.800 ;
        RECT 66.600 103.800 67.000 104.200 ;
        RECT 67.300 101.100 67.700 104.800 ;
        RECT 69.500 103.500 69.800 104.800 ;
        RECT 70.200 103.800 70.600 104.600 ;
        RECT 69.500 103.200 71.300 103.500 ;
        RECT 69.500 103.100 69.800 103.200 ;
        RECT 69.400 101.100 69.800 103.100 ;
        RECT 71.000 103.100 71.300 103.200 ;
        RECT 71.000 101.100 71.400 103.100 ;
        RECT 72.600 101.100 73.000 105.100 ;
        RECT 73.400 104.800 75.400 105.100 ;
        RECT 75.800 104.800 76.200 105.200 ;
        RECT 73.400 101.100 73.800 104.800 ;
        RECT 75.000 101.100 75.400 104.800 ;
        RECT 76.600 101.100 77.000 105.800 ;
        RECT 77.400 104.400 77.800 105.200 ;
        RECT 78.200 101.100 78.600 109.900 ;
        RECT 79.000 108.100 79.400 108.600 ;
        RECT 79.900 108.200 80.300 108.600 ;
        RECT 79.800 108.100 80.200 108.200 ;
        RECT 79.000 107.800 80.200 108.100 ;
        RECT 80.600 107.900 81.000 109.900 ;
        RECT 83.800 109.100 84.200 109.200 ;
        RECT 84.800 109.100 85.200 109.900 ;
        RECT 83.800 108.800 85.200 109.100 ;
        RECT 79.800 106.100 80.200 106.200 ;
        RECT 80.700 106.100 81.000 107.900 ;
        RECT 81.400 106.400 81.800 107.200 ;
        RECT 84.800 107.100 85.200 108.800 ;
        RECT 86.200 107.800 86.600 108.600 ;
        RECT 84.800 106.900 85.700 107.100 ;
        RECT 84.900 106.800 85.700 106.900 ;
        RECT 82.200 106.100 82.600 106.200 ;
        RECT 79.800 105.800 81.000 106.100 ;
        RECT 81.800 105.800 82.600 106.100 ;
        RECT 83.800 105.800 84.600 106.200 ;
        RECT 79.900 105.100 80.200 105.800 ;
        RECT 81.800 105.600 82.200 105.800 ;
        RECT 83.000 105.100 83.400 105.600 ;
        RECT 85.400 105.200 85.700 106.800 ;
        RECT 83.800 105.100 84.200 105.200 ;
        RECT 79.800 101.100 80.200 105.100 ;
        RECT 80.600 104.800 82.600 105.100 ;
        RECT 83.000 104.800 84.200 105.100 ;
        RECT 85.400 104.800 85.800 105.200 ;
        RECT 80.600 101.100 81.000 104.800 ;
        RECT 82.200 101.100 82.600 104.800 ;
        RECT 84.600 103.800 85.000 104.600 ;
        RECT 85.400 103.500 85.700 104.800 ;
        RECT 83.900 103.200 85.700 103.500 ;
        RECT 83.900 103.100 84.200 103.200 ;
        RECT 83.800 101.100 84.200 103.100 ;
        RECT 85.400 103.100 85.700 103.200 ;
        RECT 85.400 101.100 85.800 103.100 ;
        RECT 87.000 101.100 87.400 109.900 ;
        RECT 89.400 107.900 89.800 109.900 ;
        RECT 90.100 108.200 90.500 108.600 ;
        RECT 88.600 106.400 89.000 107.200 ;
        RECT 87.800 106.100 88.200 106.200 ;
        RECT 89.400 106.100 89.700 107.900 ;
        RECT 90.200 107.800 90.600 108.200 ;
        RECT 92.600 107.900 93.000 109.900 ;
        RECT 95.000 108.900 95.400 109.900 ;
        RECT 97.400 108.900 97.800 109.900 ;
        RECT 93.300 108.200 93.700 108.600 ;
        RECT 93.400 108.100 93.800 108.200 ;
        RECT 95.000 108.100 95.300 108.900 ;
        RECT 91.800 106.400 92.200 107.200 ;
        RECT 90.200 106.100 90.600 106.200 ;
        RECT 87.800 105.800 88.600 106.100 ;
        RECT 89.400 105.800 90.600 106.100 ;
        RECT 91.000 106.100 91.400 106.200 ;
        RECT 92.600 106.100 92.900 107.900 ;
        RECT 93.400 107.800 95.300 108.100 ;
        RECT 95.800 107.800 96.200 108.600 ;
        RECT 97.400 108.100 97.700 108.900 ;
        RECT 99.800 108.800 100.200 109.900 ;
        RECT 96.600 107.800 97.700 108.100 ;
        RECT 98.200 107.800 98.600 108.600 ;
        RECT 99.000 107.800 99.400 108.600 ;
        RECT 95.000 107.200 95.300 107.800 ;
        RECT 96.600 107.200 96.900 107.800 ;
        RECT 97.400 107.200 97.700 107.800 ;
        RECT 99.900 107.200 100.200 108.800 ;
        RECT 95.000 106.800 95.400 107.200 ;
        RECT 96.600 106.800 97.000 107.200 ;
        RECT 97.400 106.800 97.800 107.200 ;
        RECT 99.800 106.800 100.200 107.200 ;
        RECT 93.400 106.100 93.800 106.200 ;
        RECT 91.000 105.800 91.800 106.100 ;
        RECT 92.600 105.800 93.800 106.100 ;
        RECT 88.200 105.600 88.600 105.800 ;
        RECT 90.200 105.100 90.500 105.800 ;
        RECT 91.400 105.600 91.800 105.800 ;
        RECT 93.400 105.100 93.700 105.800 ;
        RECT 95.000 105.100 95.300 106.800 ;
        RECT 97.400 105.100 97.700 106.800 ;
        RECT 99.900 105.100 100.200 106.800 ;
        RECT 103.000 106.900 103.400 109.900 ;
        RECT 106.200 108.300 106.600 109.900 ;
        RECT 107.000 108.500 107.400 109.900 ;
        RECT 107.800 108.500 108.200 109.900 ;
        RECT 108.600 108.500 109.000 109.900 ;
        RECT 110.200 108.500 110.600 109.900 ;
        RECT 111.800 108.500 112.200 109.900 ;
        RECT 112.600 108.500 113.000 109.900 ;
        RECT 113.400 108.500 113.800 109.900 ;
        RECT 114.200 108.500 114.600 109.900 ;
        RECT 105.300 107.900 106.600 108.300 ;
        RECT 115.000 108.300 115.400 109.900 ;
        RECT 108.300 107.900 110.600 108.200 ;
        RECT 105.300 107.600 105.700 107.900 ;
        RECT 104.200 107.200 105.700 107.600 ;
        RECT 103.000 106.500 107.400 106.900 ;
        RECT 108.300 106.700 108.700 107.900 ;
        RECT 110.200 107.800 110.600 107.900 ;
        RECT 113.300 107.800 113.800 108.200 ;
        RECT 115.000 107.900 116.200 108.300 ;
        RECT 109.400 106.800 109.800 107.600 ;
        RECT 110.200 107.400 110.600 107.500 ;
        RECT 110.200 107.100 112.400 107.400 ;
        RECT 112.000 107.000 112.400 107.100 ;
        RECT 100.600 106.100 101.000 106.200 ;
        RECT 102.200 106.100 102.600 106.200 ;
        RECT 100.600 105.800 102.600 106.100 ;
        RECT 100.600 105.400 101.000 105.800 ;
        RECT 87.800 104.800 89.800 105.100 ;
        RECT 87.800 101.100 88.200 104.800 ;
        RECT 89.400 101.100 89.800 104.800 ;
        RECT 90.200 101.100 90.600 105.100 ;
        RECT 91.000 104.800 93.000 105.100 ;
        RECT 91.000 101.100 91.400 104.800 ;
        RECT 92.600 101.100 93.000 104.800 ;
        RECT 93.400 101.100 93.800 105.100 ;
        RECT 94.500 104.700 95.400 105.100 ;
        RECT 96.900 104.700 97.800 105.100 ;
        RECT 99.800 104.700 100.700 105.100 ;
        RECT 94.500 101.100 94.900 104.700 ;
        RECT 96.900 101.100 97.300 104.700 ;
        RECT 100.300 101.100 100.700 104.700 ;
        RECT 103.000 103.700 103.400 106.500 ;
        RECT 107.700 106.300 108.700 106.700 ;
        RECT 110.600 106.300 112.200 106.700 ;
        RECT 113.400 106.400 113.800 107.800 ;
        RECT 115.800 107.600 116.200 107.900 ;
        RECT 115.800 107.300 116.700 107.600 ;
        RECT 116.300 106.700 116.700 107.300 ;
        RECT 118.200 107.300 118.600 109.900 ;
        RECT 119.000 108.000 119.400 109.900 ;
        RECT 119.000 107.600 119.500 108.000 ;
        RECT 120.600 107.800 121.000 109.900 ;
        RECT 121.400 108.000 121.800 109.900 ;
        RECT 123.000 108.000 123.400 109.900 ;
        RECT 121.400 107.900 123.400 108.000 ;
        RECT 118.200 107.000 118.800 107.300 ;
        RECT 116.300 106.300 118.200 106.700 ;
        RECT 103.700 106.000 104.100 106.100 ;
        RECT 106.200 106.000 106.600 106.200 ;
        RECT 115.000 106.000 115.400 106.300 ;
        RECT 118.500 106.000 118.800 107.000 ;
        RECT 103.700 105.700 115.400 106.000 ;
        RECT 118.400 105.700 118.800 106.000 ;
        RECT 118.400 104.800 118.700 105.700 ;
        RECT 119.100 105.400 119.500 107.600 ;
        RECT 120.700 107.200 121.000 107.800 ;
        RECT 121.500 107.700 123.300 107.900 ;
        RECT 122.600 107.200 123.000 107.400 ;
        RECT 120.600 106.800 121.900 107.200 ;
        RECT 122.600 106.900 123.400 107.200 ;
        RECT 123.000 106.800 123.400 106.900 ;
        RECT 123.800 106.900 124.200 109.900 ;
        RECT 127.000 108.300 127.400 109.900 ;
        RECT 127.800 108.500 128.200 109.900 ;
        RECT 128.600 108.500 129.000 109.900 ;
        RECT 129.400 108.500 129.800 109.900 ;
        RECT 131.000 108.500 131.400 109.900 ;
        RECT 132.600 108.500 133.000 109.900 ;
        RECT 133.400 108.500 133.800 109.900 ;
        RECT 134.200 108.500 134.600 109.900 ;
        RECT 135.000 108.500 135.400 109.900 ;
        RECT 126.100 107.900 127.400 108.300 ;
        RECT 135.800 108.300 136.200 109.900 ;
        RECT 129.100 107.900 131.400 108.200 ;
        RECT 126.100 107.600 126.500 107.900 ;
        RECT 125.000 107.200 126.500 107.600 ;
        RECT 107.800 104.700 108.200 104.800 ;
        RECT 105.500 104.500 108.200 104.700 ;
        RECT 105.100 104.400 108.200 104.500 ;
        RECT 108.700 104.500 113.000 104.800 ;
        RECT 103.800 104.000 104.600 104.400 ;
        RECT 105.100 104.100 105.800 104.400 ;
        RECT 108.700 104.100 109.000 104.500 ;
        RECT 112.600 104.400 113.000 104.500 ;
        RECT 114.200 104.500 118.700 104.800 ;
        RECT 114.200 104.400 114.600 104.500 ;
        RECT 104.300 103.800 104.600 104.000 ;
        RECT 106.100 103.800 109.000 104.100 ;
        RECT 109.300 103.800 110.600 104.200 ;
        RECT 103.000 103.400 104.000 103.700 ;
        RECT 104.300 103.400 106.400 103.800 ;
        RECT 103.700 103.100 104.000 103.400 ;
        RECT 103.700 102.800 104.200 103.100 ;
        RECT 103.800 101.100 104.200 102.800 ;
        RECT 105.400 101.100 105.800 103.400 ;
        RECT 107.000 101.100 107.400 102.500 ;
        RECT 107.800 101.100 108.200 102.500 ;
        RECT 108.600 101.100 109.000 103.500 ;
        RECT 110.200 101.100 110.600 103.500 ;
        RECT 111.800 101.100 112.200 104.200 ;
        RECT 115.800 103.800 117.100 104.200 ;
        RECT 113.400 103.400 115.500 103.800 ;
        RECT 112.600 101.100 113.000 102.500 ;
        RECT 113.400 101.100 113.800 102.500 ;
        RECT 114.200 101.100 114.600 102.500 ;
        RECT 115.800 101.100 116.200 103.800 ;
        RECT 118.400 103.700 118.700 104.500 ;
        RECT 117.400 103.400 118.700 103.700 ;
        RECT 119.000 105.000 119.500 105.400 ;
        RECT 120.600 105.100 121.000 105.200 ;
        RECT 121.600 105.100 121.900 106.800 ;
        RECT 123.800 106.500 128.200 106.900 ;
        RECT 129.100 106.700 129.500 107.900 ;
        RECT 131.000 107.800 131.400 107.900 ;
        RECT 134.100 107.800 134.600 108.200 ;
        RECT 135.800 107.900 137.000 108.300 ;
        RECT 130.200 106.800 130.600 107.600 ;
        RECT 131.000 107.400 131.400 107.500 ;
        RECT 131.000 107.100 133.200 107.400 ;
        RECT 132.800 107.000 133.200 107.100 ;
        RECT 117.400 101.100 117.800 103.400 ;
        RECT 119.000 101.100 119.400 105.000 ;
        RECT 120.600 104.800 121.300 105.100 ;
        RECT 121.600 104.800 122.100 105.100 ;
        RECT 121.000 104.200 121.300 104.800 ;
        RECT 121.000 103.800 121.400 104.200 ;
        RECT 121.700 101.100 122.100 104.800 ;
        RECT 123.800 103.700 124.200 106.500 ;
        RECT 128.500 106.300 129.500 106.700 ;
        RECT 131.400 106.300 133.000 106.700 ;
        RECT 134.200 106.400 134.600 107.800 ;
        RECT 136.600 107.600 137.000 107.900 ;
        RECT 136.600 107.300 137.500 107.600 ;
        RECT 137.100 106.700 137.500 107.300 ;
        RECT 139.000 107.300 139.400 109.900 ;
        RECT 139.800 108.100 140.200 109.900 ;
        RECT 141.400 108.100 141.800 108.600 ;
        RECT 139.800 107.800 141.800 108.100 ;
        RECT 139.800 107.600 140.300 107.800 ;
        RECT 139.000 107.000 139.600 107.300 ;
        RECT 137.100 106.300 139.000 106.700 ;
        RECT 124.600 106.100 125.000 106.200 ;
        RECT 124.500 106.000 125.000 106.100 ;
        RECT 127.000 106.000 127.400 106.200 ;
        RECT 135.800 106.000 136.200 106.300 ;
        RECT 139.300 106.000 139.600 107.000 ;
        RECT 124.500 105.700 136.200 106.000 ;
        RECT 139.200 105.700 139.600 106.000 ;
        RECT 139.200 104.800 139.500 105.700 ;
        RECT 139.900 105.400 140.300 107.600 ;
        RECT 141.400 106.100 141.800 106.200 ;
        RECT 142.200 106.100 142.600 109.900 ;
        RECT 144.800 107.100 145.200 109.900 ;
        RECT 147.000 108.800 147.400 109.900 ;
        RECT 146.200 107.800 146.600 108.600 ;
        RECT 147.100 107.200 147.400 108.800 ;
        RECT 144.800 106.900 145.700 107.100 ;
        RECT 144.900 106.800 145.700 106.900 ;
        RECT 141.400 105.800 142.600 106.100 ;
        RECT 143.800 105.800 144.600 106.200 ;
        RECT 145.400 106.100 145.700 106.800 ;
        RECT 146.200 106.800 146.600 107.200 ;
        RECT 147.000 106.800 147.400 107.200 ;
        RECT 146.200 106.100 146.500 106.800 ;
        RECT 145.400 105.800 146.500 106.100 ;
        RECT 128.600 104.700 129.000 104.800 ;
        RECT 126.300 104.500 129.000 104.700 ;
        RECT 125.900 104.400 129.000 104.500 ;
        RECT 129.500 104.500 133.800 104.800 ;
        RECT 124.600 104.000 125.400 104.400 ;
        RECT 125.900 104.100 126.600 104.400 ;
        RECT 129.500 104.100 129.800 104.500 ;
        RECT 133.400 104.400 133.800 104.500 ;
        RECT 135.000 104.500 139.500 104.800 ;
        RECT 135.000 104.400 135.400 104.500 ;
        RECT 125.100 103.800 125.400 104.000 ;
        RECT 126.900 103.800 129.800 104.100 ;
        RECT 130.100 103.800 131.400 104.200 ;
        RECT 123.800 103.400 124.800 103.700 ;
        RECT 125.100 103.400 127.200 103.800 ;
        RECT 124.500 103.100 124.800 103.400 ;
        RECT 124.500 102.800 125.000 103.100 ;
        RECT 124.600 101.100 125.000 102.800 ;
        RECT 126.200 101.100 126.600 103.400 ;
        RECT 127.800 101.100 128.200 102.500 ;
        RECT 128.600 101.100 129.000 102.500 ;
        RECT 129.400 101.100 129.800 103.500 ;
        RECT 131.000 101.100 131.400 103.500 ;
        RECT 132.600 101.100 133.000 104.200 ;
        RECT 136.600 103.800 137.900 104.200 ;
        RECT 134.200 103.400 136.300 103.800 ;
        RECT 133.400 101.100 133.800 102.500 ;
        RECT 134.200 101.100 134.600 102.500 ;
        RECT 135.000 101.100 135.400 102.500 ;
        RECT 136.600 101.100 137.000 103.800 ;
        RECT 139.200 103.700 139.500 104.500 ;
        RECT 138.200 103.400 139.500 103.700 ;
        RECT 139.800 105.000 140.300 105.400 ;
        RECT 139.800 104.100 140.200 105.000 ;
        RECT 140.600 104.100 141.000 104.200 ;
        RECT 139.800 103.800 141.000 104.100 ;
        RECT 138.200 101.100 138.600 103.400 ;
        RECT 139.800 101.100 140.200 103.800 ;
        RECT 142.200 101.100 142.600 105.800 ;
        RECT 143.000 104.800 143.400 105.600 ;
        RECT 145.400 105.200 145.700 105.800 ;
        RECT 145.400 104.800 145.800 105.200 ;
        RECT 147.100 105.100 147.400 106.800 ;
        RECT 147.800 105.400 148.200 106.200 ;
        RECT 144.600 103.800 145.000 104.600 ;
        RECT 145.400 103.500 145.700 104.800 ;
        RECT 147.000 104.700 147.900 105.100 ;
        RECT 143.900 103.200 145.700 103.500 ;
        RECT 143.900 103.100 144.200 103.200 ;
        RECT 143.800 101.100 144.200 103.100 ;
        RECT 145.400 103.100 145.700 103.200 ;
        RECT 145.400 101.100 145.800 103.100 ;
        RECT 147.500 101.100 147.900 104.700 ;
        RECT 0.600 97.900 1.000 99.900 ;
        RECT 0.700 97.800 1.000 97.900 ;
        RECT 2.200 97.900 2.600 99.900 ;
        RECT 2.200 97.800 2.500 97.900 ;
        RECT 0.700 97.500 2.500 97.800 ;
        RECT 0.700 96.200 1.000 97.500 ;
        RECT 1.400 96.400 1.800 97.200 ;
        RECT 0.600 95.800 1.000 96.200 ;
        RECT 0.700 94.200 1.000 95.800 ;
        RECT 3.000 95.400 3.400 96.200 ;
        RECT 1.400 94.800 2.600 95.200 ;
        RECT 0.700 94.100 1.500 94.200 ;
        RECT 0.700 93.900 1.600 94.100 ;
        RECT 1.200 91.100 1.600 93.900 ;
        RECT 3.800 93.400 4.200 94.200 ;
        RECT 4.600 91.100 5.000 99.900 ;
        RECT 5.400 97.900 5.800 99.900 ;
        RECT 5.500 97.800 5.800 97.900 ;
        RECT 7.000 97.900 7.400 99.900 ;
        RECT 7.000 97.800 7.300 97.900 ;
        RECT 5.500 97.500 7.300 97.800 ;
        RECT 5.500 96.200 5.800 97.500 ;
        RECT 6.200 96.400 6.600 97.200 ;
        RECT 5.400 95.800 5.800 96.200 ;
        RECT 5.500 94.200 5.800 95.800 ;
        RECT 7.800 95.400 8.200 96.200 ;
        RECT 8.600 96.100 9.000 96.200 ;
        RECT 9.400 96.100 9.800 99.900 ;
        RECT 8.600 95.800 9.800 96.100 ;
        RECT 6.600 94.800 7.400 95.200 ;
        RECT 5.500 94.100 6.300 94.200 ;
        RECT 5.500 93.900 6.400 94.100 ;
        RECT 6.000 91.100 6.400 93.900 ;
        RECT 8.600 93.400 9.000 94.200 ;
        RECT 9.400 93.100 9.800 95.800 ;
        RECT 10.200 95.800 10.600 96.600 ;
        RECT 11.000 96.200 11.400 99.900 ;
        RECT 12.600 99.600 14.600 99.900 ;
        RECT 12.600 96.200 13.000 99.600 ;
        RECT 11.000 95.900 13.000 96.200 ;
        RECT 13.400 95.900 13.800 99.300 ;
        RECT 14.200 95.900 14.600 99.600 ;
        RECT 15.000 97.900 15.400 99.900 ;
        RECT 15.100 97.800 15.400 97.900 ;
        RECT 16.600 97.900 17.000 99.900 ;
        RECT 16.600 97.800 16.900 97.900 ;
        RECT 15.100 97.500 16.900 97.800 ;
        RECT 15.100 96.200 15.400 97.500 ;
        RECT 15.800 96.400 16.200 97.200 ;
        RECT 18.200 96.200 18.600 99.900 ;
        RECT 19.800 96.200 20.200 99.900 ;
        RECT 10.200 95.100 10.500 95.800 ;
        RECT 13.400 95.600 13.700 95.900 ;
        RECT 15.000 95.800 15.400 96.200 ;
        RECT 11.400 95.200 11.800 95.400 ;
        RECT 12.700 95.300 13.700 95.600 ;
        RECT 12.700 95.200 13.000 95.300 ;
        RECT 11.000 95.100 11.800 95.200 ;
        RECT 10.200 94.900 11.800 95.100 ;
        RECT 10.200 94.800 11.400 94.900 ;
        RECT 12.600 94.800 13.000 95.200 ;
        RECT 14.200 94.800 14.600 95.600 ;
        RECT 11.800 93.800 12.200 94.600 ;
        RECT 12.700 94.200 13.000 94.800 ;
        RECT 13.300 94.400 13.700 94.800 ;
        RECT 12.600 93.800 13.000 94.200 ;
        RECT 13.400 94.200 13.700 94.400 ;
        RECT 15.100 94.200 15.400 95.800 ;
        RECT 17.400 95.400 17.800 96.200 ;
        RECT 18.200 95.900 20.200 96.200 ;
        RECT 20.600 95.900 21.000 99.900 ;
        RECT 22.700 99.200 23.100 99.900 ;
        RECT 22.200 98.800 23.100 99.200 ;
        RECT 22.700 96.200 23.100 98.800 ;
        RECT 23.400 96.800 23.800 97.200 ;
        RECT 23.500 96.200 23.800 96.800 ;
        RECT 22.700 95.900 23.200 96.200 ;
        RECT 23.500 95.900 24.200 96.200 ;
        RECT 24.600 95.900 25.000 99.900 ;
        RECT 25.400 96.200 25.800 99.900 ;
        RECT 27.000 96.200 27.400 99.900 ;
        RECT 27.800 97.900 28.200 99.900 ;
        RECT 27.900 97.800 28.200 97.900 ;
        RECT 29.400 97.900 29.800 99.900 ;
        RECT 31.000 97.900 31.400 99.900 ;
        RECT 29.400 97.800 29.700 97.900 ;
        RECT 27.900 97.500 29.700 97.800 ;
        RECT 31.100 97.800 31.400 97.900 ;
        RECT 32.600 97.900 33.000 99.900 ;
        RECT 32.600 97.800 32.900 97.900 ;
        RECT 31.100 97.500 32.900 97.800 ;
        RECT 27.900 96.200 28.200 97.500 ;
        RECT 28.600 96.400 29.000 97.200 ;
        RECT 31.100 96.200 31.400 97.500 ;
        RECT 31.800 96.400 32.200 97.200 ;
        RECT 25.400 95.900 27.400 96.200 ;
        RECT 18.600 95.200 19.000 95.400 ;
        RECT 20.600 95.200 20.900 95.900 ;
        RECT 16.200 94.800 17.000 95.200 ;
        RECT 18.200 94.900 19.000 95.200 ;
        RECT 19.800 94.900 21.000 95.200 ;
        RECT 18.200 94.800 18.600 94.900 ;
        RECT 13.400 93.800 13.800 94.200 ;
        RECT 15.100 94.100 15.900 94.200 ;
        RECT 15.100 93.900 16.000 94.100 ;
        RECT 12.700 93.100 13.000 93.800 ;
        RECT 9.400 92.800 10.300 93.100 ;
        RECT 9.900 91.100 10.300 92.800 ;
        RECT 12.500 91.100 13.300 93.100 ;
        RECT 15.600 91.100 16.000 93.900 ;
        RECT 19.000 93.800 19.400 94.600 ;
        RECT 19.800 94.100 20.100 94.900 ;
        RECT 20.600 94.800 21.000 94.900 ;
        RECT 22.200 94.400 22.600 95.200 ;
        RECT 22.900 94.200 23.200 95.900 ;
        RECT 23.800 95.800 24.200 95.900 ;
        RECT 24.700 95.200 25.000 95.900 ;
        RECT 27.800 95.800 28.200 96.200 ;
        RECT 26.600 95.200 27.000 95.400 ;
        RECT 24.600 94.900 25.800 95.200 ;
        RECT 26.600 94.900 27.400 95.200 ;
        RECT 24.600 94.800 25.000 94.900 ;
        RECT 21.400 94.100 21.800 94.200 ;
        RECT 19.800 93.800 22.200 94.100 ;
        RECT 22.900 93.800 24.200 94.200 ;
        RECT 19.800 93.100 20.100 93.800 ;
        RECT 21.800 93.600 22.200 93.800 ;
        RECT 19.800 91.100 20.200 93.100 ;
        RECT 20.600 92.800 21.000 93.200 ;
        RECT 21.500 93.100 23.300 93.300 ;
        RECT 23.800 93.100 24.100 93.800 ;
        RECT 21.400 93.000 23.400 93.100 ;
        RECT 20.500 92.400 20.900 92.800 ;
        RECT 21.400 91.100 21.800 93.000 ;
        RECT 23.000 91.100 23.400 93.000 ;
        RECT 23.800 91.100 24.200 93.100 ;
        RECT 24.600 92.800 25.000 93.200 ;
        RECT 25.500 93.100 25.800 94.900 ;
        RECT 27.000 94.800 27.400 94.900 ;
        RECT 26.200 93.800 26.600 94.600 ;
        RECT 27.900 94.200 28.200 95.800 ;
        RECT 30.200 95.400 30.600 96.200 ;
        RECT 31.000 95.800 31.400 96.200 ;
        RECT 29.000 94.800 29.800 95.200 ;
        RECT 31.100 94.200 31.400 95.800 ;
        RECT 33.400 95.400 33.800 96.200 ;
        RECT 34.200 95.900 34.600 99.900 ;
        RECT 35.000 96.200 35.400 99.900 ;
        RECT 36.600 96.200 37.000 99.900 ;
        RECT 38.200 97.800 38.600 99.900 ;
        RECT 39.800 97.900 40.200 99.900 ;
        RECT 39.800 97.800 40.100 97.900 ;
        RECT 38.200 97.500 40.100 97.800 ;
        RECT 38.200 97.200 38.500 97.500 ;
        RECT 38.200 96.800 38.600 97.200 ;
        RECT 39.000 96.400 39.400 97.200 ;
        RECT 39.800 96.200 40.100 97.500 ;
        RECT 35.000 95.900 37.000 96.200 ;
        RECT 34.300 95.200 34.600 95.900 ;
        RECT 37.400 95.400 37.800 96.200 ;
        RECT 39.800 95.800 40.200 96.200 ;
        RECT 36.200 95.200 36.600 95.400 ;
        RECT 32.200 94.800 33.000 95.200 ;
        RECT 34.200 94.900 35.400 95.200 ;
        RECT 36.200 94.900 37.000 95.200 ;
        RECT 34.200 94.800 34.600 94.900 ;
        RECT 35.100 94.200 35.400 94.900 ;
        RECT 36.600 94.800 37.000 94.900 ;
        RECT 38.200 94.800 39.000 95.200 ;
        RECT 27.900 94.100 28.700 94.200 ;
        RECT 31.100 94.100 31.900 94.200 ;
        RECT 27.900 93.900 28.800 94.100 ;
        RECT 31.100 93.900 32.000 94.100 ;
        RECT 24.700 92.400 25.100 92.800 ;
        RECT 25.400 91.100 25.800 93.100 ;
        RECT 28.400 91.100 28.800 93.900 ;
        RECT 31.600 91.100 32.000 93.900 ;
        RECT 35.000 93.800 35.400 94.200 ;
        RECT 35.800 93.800 36.200 94.600 ;
        RECT 39.800 94.200 40.100 95.800 ;
        RECT 39.300 94.100 40.100 94.200 ;
        RECT 39.200 93.900 40.100 94.100 ;
        RECT 34.200 92.800 34.600 93.200 ;
        RECT 35.100 93.100 35.400 93.800 ;
        RECT 34.300 92.400 34.700 92.800 ;
        RECT 35.000 91.100 35.400 93.100 ;
        RECT 39.200 91.100 39.600 93.900 ;
        RECT 40.600 91.100 41.000 99.900 ;
        RECT 43.000 97.900 43.400 99.900 ;
        RECT 43.100 97.800 43.400 97.900 ;
        RECT 44.600 97.900 45.000 99.900 ;
        RECT 46.200 97.900 46.600 99.900 ;
        RECT 44.600 97.800 44.900 97.900 ;
        RECT 43.100 97.500 44.900 97.800 ;
        RECT 46.300 97.800 46.600 97.900 ;
        RECT 47.800 97.900 48.200 99.900 ;
        RECT 51.000 97.900 51.400 99.900 ;
        RECT 47.800 97.800 48.100 97.900 ;
        RECT 46.300 97.500 48.100 97.800 ;
        RECT 51.100 97.800 51.400 97.900 ;
        RECT 52.600 97.900 53.000 99.900 ;
        RECT 52.600 97.800 52.900 97.900 ;
        RECT 54.200 97.800 54.600 99.900 ;
        RECT 55.800 97.900 56.200 99.900 ;
        RECT 56.900 99.200 57.300 99.900 ;
        RECT 56.600 98.800 57.300 99.200 ;
        RECT 55.800 97.800 56.100 97.900 ;
        RECT 51.100 97.500 52.900 97.800 ;
        RECT 54.300 97.500 56.100 97.800 ;
        RECT 43.800 96.400 44.200 97.200 ;
        RECT 44.600 97.100 44.900 97.500 ;
        RECT 47.000 97.100 47.400 97.200 ;
        RECT 44.600 96.800 47.400 97.100 ;
        RECT 44.600 96.200 44.900 96.800 ;
        RECT 47.000 96.400 47.400 96.800 ;
        RECT 47.800 96.200 48.100 97.500 ;
        RECT 51.800 96.400 52.200 97.200 ;
        RECT 52.600 96.200 52.900 97.500 ;
        RECT 55.000 96.400 55.400 97.200 ;
        RECT 55.800 96.200 56.100 97.500 ;
        RECT 56.900 96.300 57.300 98.800 ;
        RECT 59.000 97.900 59.400 99.900 ;
        RECT 59.100 97.800 59.400 97.900 ;
        RECT 60.600 97.900 61.000 99.900 ;
        RECT 60.600 97.800 60.900 97.900 ;
        RECT 59.100 97.500 60.900 97.800 ;
        RECT 42.200 95.400 42.600 96.200 ;
        RECT 44.600 95.800 45.000 96.200 ;
        RECT 43.000 94.800 43.800 95.200 ;
        RECT 44.600 94.200 44.900 95.800 ;
        RECT 45.400 95.400 45.800 96.200 ;
        RECT 47.800 95.800 48.200 96.200 ;
        RECT 46.200 94.800 47.000 95.200 ;
        RECT 47.800 94.200 48.100 95.800 ;
        RECT 50.200 95.400 50.600 96.200 ;
        RECT 52.600 95.800 53.000 96.200 ;
        RECT 51.000 94.800 51.800 95.200 ;
        RECT 52.600 94.200 52.900 95.800 ;
        RECT 53.400 95.400 53.800 96.200 ;
        RECT 55.800 95.800 56.200 96.200 ;
        RECT 56.900 95.900 57.800 96.300 ;
        RECT 59.100 96.200 59.400 97.500 ;
        RECT 59.800 96.400 60.200 97.200 ;
        RECT 54.200 94.800 55.000 95.200 ;
        RECT 55.800 94.200 56.100 95.800 ;
        RECT 56.600 94.800 57.000 95.600 ;
        RECT 41.400 93.400 41.800 94.200 ;
        RECT 44.100 94.100 44.900 94.200 ;
        RECT 47.300 94.100 48.100 94.200 ;
        RECT 52.100 94.100 52.900 94.200 ;
        RECT 55.300 94.100 56.100 94.200 ;
        RECT 44.000 93.900 44.900 94.100 ;
        RECT 47.200 93.900 48.100 94.100 ;
        RECT 52.000 93.900 52.900 94.100 ;
        RECT 55.200 93.900 56.100 94.100 ;
        RECT 57.400 94.200 57.700 95.900 ;
        RECT 59.000 95.800 59.400 96.200 ;
        RECT 59.100 94.200 59.400 95.800 ;
        RECT 61.400 95.400 61.800 96.200 ;
        RECT 62.200 95.900 62.600 99.900 ;
        RECT 63.000 96.200 63.400 99.900 ;
        RECT 64.600 96.200 65.000 99.900 ;
        RECT 63.000 95.900 65.000 96.200 ;
        RECT 65.400 95.900 65.800 99.900 ;
        RECT 66.200 96.200 66.600 99.900 ;
        RECT 67.800 96.200 68.200 99.900 ;
        RECT 69.400 97.900 69.800 99.900 ;
        RECT 69.500 97.800 69.800 97.900 ;
        RECT 71.000 97.900 71.400 99.900 ;
        RECT 71.000 97.800 71.300 97.900 ;
        RECT 69.500 97.500 71.300 97.800 ;
        RECT 70.200 96.400 70.600 97.200 ;
        RECT 71.000 96.200 71.300 97.500 ;
        RECT 66.200 95.900 68.200 96.200 ;
        RECT 62.300 95.200 62.600 95.900 ;
        RECT 64.200 95.200 64.600 95.400 ;
        RECT 65.500 95.200 65.800 95.900 ;
        RECT 68.600 95.400 69.000 96.200 ;
        RECT 71.000 95.800 71.400 96.200 ;
        RECT 71.800 95.900 72.200 99.900 ;
        RECT 72.600 96.200 73.000 99.900 ;
        RECT 74.200 96.200 74.600 99.900 ;
        RECT 72.600 95.900 74.600 96.200 ;
        RECT 75.300 96.300 75.700 99.900 ;
        RECT 78.700 97.200 79.700 99.900 ;
        RECT 82.500 99.200 82.900 99.900 ;
        RECT 85.900 99.200 86.300 99.900 ;
        RECT 82.500 98.800 83.400 99.200 ;
        RECT 85.400 98.800 86.300 99.200 ;
        RECT 78.200 96.800 79.700 97.200 ;
        RECT 75.300 95.900 76.200 96.300 ;
        RECT 78.700 95.900 79.700 96.800 ;
        RECT 81.800 96.800 82.200 97.200 ;
        RECT 81.800 96.200 82.100 96.800 ;
        RECT 82.500 96.200 82.900 98.800 ;
        RECT 81.400 95.900 82.100 96.200 ;
        RECT 82.400 95.900 82.900 96.200 ;
        RECT 85.900 96.200 86.300 98.800 ;
        RECT 86.600 96.800 87.000 97.200 ;
        RECT 86.700 96.200 87.000 96.800 ;
        RECT 85.900 95.900 86.400 96.200 ;
        RECT 86.700 96.100 87.400 96.200 ;
        RECT 87.800 96.100 88.200 99.900 ;
        RECT 90.500 99.200 90.900 99.900 ;
        RECT 90.500 98.800 91.400 99.200 ;
        RECT 89.800 96.800 90.200 97.200 ;
        RECT 89.800 96.200 90.100 96.800 ;
        RECT 90.500 96.200 90.900 98.800 ;
        RECT 86.700 95.900 88.200 96.100 ;
        RECT 67.400 95.200 67.800 95.400 ;
        RECT 60.200 94.800 61.000 95.200 ;
        RECT 62.200 94.900 63.400 95.200 ;
        RECT 64.200 94.900 65.000 95.200 ;
        RECT 62.200 94.800 62.600 94.900 ;
        RECT 44.000 91.100 44.400 93.900 ;
        RECT 47.200 91.100 47.600 93.900 ;
        RECT 52.000 91.100 52.400 93.900 ;
        RECT 55.200 91.100 55.600 93.900 ;
        RECT 57.400 93.800 57.800 94.200 ;
        RECT 59.100 94.100 59.900 94.200 ;
        RECT 59.100 93.900 60.000 94.100 ;
        RECT 57.400 92.100 57.700 93.800 ;
        RECT 58.200 92.400 58.600 93.200 ;
        RECT 57.400 91.100 57.800 92.100 ;
        RECT 59.600 91.100 60.000 93.900 ;
        RECT 62.200 92.800 62.600 93.200 ;
        RECT 63.100 93.100 63.400 94.900 ;
        RECT 64.600 94.800 65.000 94.900 ;
        RECT 65.400 94.900 66.600 95.200 ;
        RECT 67.400 94.900 68.200 95.200 ;
        RECT 65.400 94.800 65.800 94.900 ;
        RECT 63.800 93.800 64.200 94.600 ;
        RECT 62.300 92.400 62.700 92.800 ;
        RECT 63.000 91.100 63.400 93.100 ;
        RECT 65.400 92.800 65.800 93.200 ;
        RECT 66.300 93.100 66.600 94.900 ;
        RECT 67.800 94.800 68.200 94.900 ;
        RECT 69.400 94.800 70.200 95.200 ;
        RECT 67.000 94.100 67.400 94.600 ;
        RECT 71.000 94.200 71.300 95.800 ;
        RECT 71.900 95.200 72.200 95.900 ;
        RECT 73.800 95.200 74.200 95.400 ;
        RECT 67.800 94.100 68.200 94.200 ;
        RECT 70.500 94.100 71.300 94.200 ;
        RECT 67.000 93.800 68.200 94.100 ;
        RECT 70.400 93.900 71.300 94.100 ;
        RECT 71.800 94.900 73.000 95.200 ;
        RECT 73.800 94.900 74.600 95.200 ;
        RECT 71.800 94.800 72.200 94.900 ;
        RECT 71.800 94.200 72.100 94.800 ;
        RECT 65.500 92.400 65.900 92.800 ;
        RECT 66.200 91.100 66.600 93.100 ;
        RECT 70.400 91.100 70.800 93.900 ;
        RECT 71.800 93.800 72.200 94.200 ;
        RECT 71.800 92.800 72.200 93.200 ;
        RECT 72.700 93.100 73.000 94.900 ;
        RECT 74.200 94.800 74.600 94.900 ;
        RECT 75.000 94.800 75.400 95.600 ;
        RECT 73.400 93.800 73.800 94.600 ;
        RECT 75.800 94.200 76.100 95.900 ;
        RECT 76.600 95.100 77.000 95.200 ;
        RECT 78.200 95.100 78.600 95.200 ;
        RECT 76.600 94.800 78.600 95.100 ;
        RECT 78.200 94.400 78.600 94.800 ;
        RECT 79.000 94.200 79.300 95.900 ;
        RECT 81.400 95.800 81.800 95.900 ;
        RECT 79.800 94.400 80.200 95.200 ;
        RECT 75.000 93.800 75.400 94.200 ;
        RECT 75.800 93.800 76.200 94.200 ;
        RECT 77.400 94.100 77.800 94.200 ;
        RECT 79.000 94.100 79.400 94.200 ;
        RECT 76.600 93.800 78.200 94.100 ;
        RECT 79.000 93.800 80.200 94.100 ;
        RECT 80.600 93.800 81.000 94.600 ;
        RECT 82.400 94.200 82.700 95.900 ;
        RECT 83.000 95.100 83.400 95.200 ;
        RECT 85.400 95.100 85.800 95.200 ;
        RECT 83.000 94.800 85.800 95.100 ;
        RECT 83.000 94.400 83.400 94.800 ;
        RECT 85.400 94.400 85.800 94.800 ;
        RECT 86.100 94.200 86.400 95.900 ;
        RECT 87.000 95.800 88.200 95.900 ;
        RECT 89.400 95.900 90.100 96.200 ;
        RECT 90.400 95.900 90.900 96.200 ;
        RECT 92.900 96.300 93.300 99.900 ;
        RECT 95.000 97.900 95.400 99.900 ;
        RECT 95.100 97.800 95.400 97.900 ;
        RECT 96.600 97.900 97.000 99.900 ;
        RECT 96.600 97.800 96.900 97.900 ;
        RECT 95.100 97.500 96.900 97.800 ;
        RECT 92.900 95.900 93.800 96.300 ;
        RECT 95.100 96.200 95.400 97.500 ;
        RECT 96.600 97.200 96.900 97.500 ;
        RECT 95.800 96.400 96.200 97.200 ;
        RECT 96.600 96.800 97.000 97.200 ;
        RECT 99.500 96.200 99.900 99.900 ;
        RECT 100.200 96.800 100.600 97.200 ;
        RECT 100.300 96.200 100.600 96.800 ;
        RECT 104.300 96.200 104.700 99.900 ;
        RECT 105.000 96.800 105.400 97.200 ;
        RECT 105.100 96.200 105.400 96.800 ;
        RECT 89.400 95.800 89.800 95.900 ;
        RECT 87.000 95.200 87.300 95.800 ;
        RECT 87.000 94.800 87.400 95.200 ;
        RECT 81.400 93.800 82.700 94.200 ;
        RECT 83.800 94.100 84.200 94.200 ;
        RECT 84.600 94.100 85.000 94.200 ;
        RECT 83.400 93.800 85.400 94.100 ;
        RECT 86.100 93.800 87.400 94.200 ;
        RECT 71.900 92.400 72.300 92.800 ;
        RECT 72.600 91.100 73.000 93.100 ;
        RECT 75.000 93.100 75.300 93.800 ;
        RECT 75.800 93.100 76.100 93.800 ;
        RECT 75.000 92.800 76.100 93.100 ;
        RECT 75.800 92.100 76.100 92.800 ;
        RECT 76.600 93.200 76.900 93.800 ;
        RECT 77.800 93.600 78.200 93.800 ;
        RECT 76.600 92.400 77.000 93.200 ;
        RECT 77.500 93.100 79.300 93.300 ;
        RECT 79.900 93.100 80.200 93.800 ;
        RECT 81.500 93.100 81.800 93.800 ;
        RECT 83.400 93.600 83.800 93.800 ;
        RECT 85.000 93.600 85.400 93.800 ;
        RECT 82.300 93.100 84.100 93.300 ;
        RECT 84.700 93.100 86.500 93.300 ;
        RECT 87.000 93.100 87.300 93.800 ;
        RECT 77.400 93.000 79.400 93.100 ;
        RECT 75.800 91.100 76.200 92.100 ;
        RECT 77.400 91.100 77.800 93.000 ;
        RECT 79.000 91.400 79.400 93.000 ;
        RECT 79.800 91.700 80.200 93.100 ;
        RECT 80.600 91.400 81.000 93.100 ;
        RECT 79.000 91.100 81.000 91.400 ;
        RECT 81.400 91.100 81.800 93.100 ;
        RECT 82.200 93.000 84.200 93.100 ;
        RECT 82.200 91.100 82.600 93.000 ;
        RECT 83.800 91.100 84.200 93.000 ;
        RECT 84.600 93.000 86.600 93.100 ;
        RECT 84.600 91.100 85.000 93.000 ;
        RECT 86.200 91.100 86.600 93.000 ;
        RECT 87.000 91.100 87.400 93.100 ;
        RECT 87.800 91.100 88.200 95.800 ;
        RECT 90.400 94.200 90.700 95.900 ;
        RECT 91.000 94.400 91.400 95.200 ;
        RECT 92.600 94.800 93.000 95.600 ;
        RECT 93.400 94.200 93.700 95.900 ;
        RECT 95.000 95.800 95.400 96.200 ;
        RECT 95.100 94.200 95.400 95.800 ;
        RECT 97.400 95.400 97.800 96.200 ;
        RECT 99.000 95.800 100.000 96.200 ;
        RECT 100.300 96.100 101.000 96.200 ;
        RECT 102.200 96.100 102.600 96.200 ;
        RECT 100.300 95.900 102.600 96.100 ;
        RECT 104.300 95.900 104.800 96.200 ;
        RECT 105.100 95.900 105.800 96.200 ;
        RECT 100.600 95.800 102.600 95.900 ;
        RECT 96.200 94.800 97.000 95.200 ;
        RECT 99.000 94.400 99.400 95.200 ;
        RECT 99.700 94.200 100.000 95.800 ;
        RECT 103.800 94.400 104.200 95.200 ;
        RECT 104.500 94.200 104.800 95.900 ;
        RECT 105.400 95.800 105.800 95.900 ;
        RECT 105.400 94.800 105.800 95.200 ;
        RECT 105.400 94.200 105.700 94.800 ;
        RECT 88.600 93.400 89.000 94.200 ;
        RECT 89.400 93.800 90.700 94.200 ;
        RECT 91.800 94.100 92.200 94.200 ;
        RECT 91.400 93.800 92.200 94.100 ;
        RECT 93.400 93.800 93.800 94.200 ;
        RECT 95.100 94.100 95.900 94.200 ;
        RECT 98.200 94.100 98.600 94.200 ;
        RECT 95.100 93.900 96.000 94.100 ;
        RECT 89.500 93.100 89.800 93.800 ;
        RECT 91.400 93.600 91.800 93.800 ;
        RECT 90.300 93.100 92.100 93.300 ;
        RECT 92.600 93.100 93.000 93.200 ;
        RECT 93.400 93.100 93.700 93.800 ;
        RECT 89.400 91.100 89.800 93.100 ;
        RECT 90.200 93.000 92.200 93.100 ;
        RECT 90.200 91.100 90.600 93.000 ;
        RECT 91.800 91.100 92.200 93.000 ;
        RECT 92.600 92.800 93.700 93.100 ;
        RECT 93.400 92.100 93.700 92.800 ;
        RECT 94.200 92.400 94.600 93.200 ;
        RECT 93.400 91.100 93.800 92.100 ;
        RECT 95.600 91.100 96.000 93.900 ;
        RECT 98.200 93.800 99.000 94.100 ;
        RECT 99.700 93.800 101.000 94.200 ;
        RECT 103.000 94.100 103.400 94.200 ;
        RECT 103.000 93.800 103.800 94.100 ;
        RECT 104.500 93.800 105.800 94.200 ;
        RECT 98.600 93.600 99.000 93.800 ;
        RECT 98.300 93.100 100.100 93.300 ;
        RECT 100.600 93.100 100.900 93.800 ;
        RECT 103.400 93.600 103.800 93.800 ;
        RECT 103.100 93.100 104.900 93.300 ;
        RECT 105.400 93.100 105.700 93.800 ;
        RECT 98.200 93.000 100.200 93.100 ;
        RECT 98.200 91.100 98.600 93.000 ;
        RECT 99.800 91.100 100.200 93.000 ;
        RECT 100.600 91.100 101.000 93.100 ;
        RECT 103.000 93.000 105.000 93.100 ;
        RECT 103.000 91.100 103.400 93.000 ;
        RECT 104.600 91.100 105.000 93.000 ;
        RECT 105.400 91.100 105.800 93.100 ;
        RECT 106.200 91.100 106.600 99.900 ;
        RECT 108.100 96.300 108.500 99.900 ;
        RECT 110.500 96.300 110.900 99.900 ;
        RECT 108.100 95.900 109.000 96.300 ;
        RECT 110.500 95.900 111.400 96.300 ;
        RECT 107.800 94.800 108.200 95.600 ;
        RECT 108.600 94.200 108.900 95.900 ;
        RECT 110.200 94.800 110.600 95.600 ;
        RECT 111.000 95.100 111.300 95.900 ;
        RECT 112.600 95.800 113.000 96.600 ;
        RECT 112.600 95.100 112.900 95.800 ;
        RECT 111.000 94.800 112.900 95.100 ;
        RECT 113.400 95.100 113.800 99.900 ;
        RECT 116.300 99.200 116.700 99.900 ;
        RECT 115.800 98.800 116.700 99.200 ;
        RECT 116.300 96.200 116.700 98.800 ;
        RECT 118.200 96.200 118.600 99.900 ;
        RECT 119.800 96.200 120.200 99.900 ;
        RECT 116.300 95.900 116.800 96.200 ;
        RECT 118.200 95.900 120.200 96.200 ;
        RECT 120.600 95.900 121.000 99.900 ;
        RECT 122.700 96.300 123.100 99.900 ;
        RECT 124.600 98.200 125.000 99.900 ;
        RECT 124.500 97.900 125.000 98.200 ;
        RECT 124.500 97.600 124.800 97.900 ;
        RECT 126.200 97.600 126.600 99.900 ;
        RECT 127.800 98.500 128.200 99.900 ;
        RECT 128.600 98.500 129.000 99.900 ;
        RECT 122.200 95.900 123.100 96.300 ;
        RECT 123.800 97.300 124.800 97.600 ;
        RECT 113.400 94.800 115.300 95.100 ;
        RECT 111.000 94.200 111.300 94.800 ;
        RECT 108.600 93.800 109.000 94.200 ;
        RECT 111.000 93.800 111.400 94.200 ;
        RECT 107.000 93.100 107.400 93.200 ;
        RECT 108.600 93.100 108.900 93.800 ;
        RECT 107.000 92.800 108.900 93.100 ;
        RECT 107.000 92.400 107.400 92.800 ;
        RECT 108.600 92.100 108.900 92.800 ;
        RECT 109.400 92.400 109.800 93.200 ;
        RECT 111.000 92.100 111.300 93.800 ;
        RECT 111.800 92.400 112.200 93.200 ;
        RECT 113.400 93.100 113.800 94.800 ;
        RECT 115.000 94.200 115.300 94.800 ;
        RECT 115.800 94.400 116.200 95.200 ;
        RECT 116.500 94.200 116.800 95.900 ;
        RECT 118.600 95.200 119.000 95.400 ;
        RECT 120.600 95.200 120.900 95.900 ;
        RECT 118.200 94.900 119.000 95.200 ;
        RECT 119.800 94.900 121.000 95.200 ;
        RECT 118.200 94.800 118.600 94.900 ;
        RECT 114.200 93.400 114.600 94.200 ;
        RECT 115.000 94.100 115.400 94.200 ;
        RECT 115.000 93.800 115.800 94.100 ;
        RECT 116.500 93.800 117.800 94.200 ;
        RECT 119.000 93.800 119.400 94.600 ;
        RECT 115.400 93.600 115.800 93.800 ;
        RECT 115.100 93.100 116.900 93.300 ;
        RECT 117.400 93.100 117.700 93.800 ;
        RECT 119.800 93.100 120.100 94.900 ;
        RECT 120.600 94.800 121.000 94.900 ;
        RECT 122.300 94.200 122.600 95.900 ;
        RECT 122.200 94.100 122.600 94.200 ;
        RECT 120.600 93.800 122.600 94.100 ;
        RECT 120.600 93.200 120.900 93.800 ;
        RECT 112.900 92.800 113.800 93.100 ;
        RECT 115.000 93.000 117.000 93.100 ;
        RECT 108.600 91.100 109.000 92.100 ;
        RECT 111.000 91.100 111.400 92.100 ;
        RECT 112.900 91.100 113.300 92.800 ;
        RECT 115.000 91.100 115.400 93.000 ;
        RECT 116.600 91.100 117.000 93.000 ;
        RECT 117.400 91.100 117.800 93.100 ;
        RECT 119.800 91.100 120.200 93.100 ;
        RECT 120.600 92.800 121.000 93.200 ;
        RECT 120.500 92.400 120.900 92.800 ;
        RECT 121.400 92.400 121.800 93.200 ;
        RECT 122.300 92.100 122.600 93.800 ;
        RECT 122.200 91.100 122.600 92.100 ;
        RECT 123.800 94.500 124.200 97.300 ;
        RECT 125.100 97.200 127.200 97.600 ;
        RECT 129.400 97.500 129.800 99.900 ;
        RECT 131.000 97.500 131.400 99.900 ;
        RECT 125.100 97.000 125.400 97.200 ;
        RECT 124.600 96.600 125.400 97.000 ;
        RECT 126.900 96.900 129.800 97.200 ;
        RECT 125.900 96.600 126.600 96.900 ;
        RECT 125.900 96.500 129.000 96.600 ;
        RECT 126.300 96.300 129.000 96.500 ;
        RECT 128.600 96.200 129.000 96.300 ;
        RECT 129.500 96.500 129.800 96.900 ;
        RECT 130.100 96.800 131.400 97.200 ;
        RECT 132.600 96.800 133.000 99.900 ;
        RECT 133.400 98.500 133.800 99.900 ;
        RECT 134.200 98.500 134.600 99.900 ;
        RECT 135.000 98.500 135.400 99.900 ;
        RECT 134.200 97.200 136.300 97.600 ;
        RECT 136.600 97.200 137.000 99.900 ;
        RECT 138.200 97.600 138.600 99.900 ;
        RECT 138.200 97.300 139.500 97.600 ;
        RECT 136.600 96.800 137.900 97.200 ;
        RECT 133.400 96.500 133.800 96.600 ;
        RECT 129.500 96.200 133.800 96.500 ;
        RECT 135.000 96.500 135.400 96.600 ;
        RECT 139.200 96.500 139.500 97.300 ;
        RECT 135.000 96.200 139.500 96.500 ;
        RECT 139.200 95.300 139.500 96.200 ;
        RECT 139.800 96.000 140.200 99.900 ;
        RECT 141.400 96.200 141.800 99.900 ;
        RECT 145.100 99.200 145.500 99.900 ;
        RECT 144.600 98.800 145.500 99.200 ;
        RECT 145.100 96.300 145.500 98.800 ;
        RECT 139.800 95.600 140.300 96.000 ;
        RECT 141.400 95.900 142.500 96.200 ;
        RECT 144.600 95.900 145.500 96.300 ;
        RECT 146.200 96.200 146.600 99.900 ;
        RECT 146.200 95.900 147.300 96.200 ;
        RECT 124.500 95.000 136.200 95.300 ;
        RECT 139.200 95.000 139.600 95.300 ;
        RECT 124.500 94.900 124.900 95.000 ;
        RECT 127.000 94.800 127.400 95.000 ;
        RECT 135.800 94.700 136.200 95.000 ;
        RECT 123.800 94.100 128.200 94.500 ;
        RECT 128.500 94.300 129.500 94.700 ;
        RECT 131.400 94.300 133.000 94.700 ;
        RECT 123.800 91.100 124.200 94.100 ;
        RECT 125.000 93.400 126.500 93.800 ;
        RECT 126.100 93.100 126.500 93.400 ;
        RECT 129.100 93.100 129.500 94.300 ;
        RECT 130.200 93.400 130.600 94.200 ;
        RECT 132.800 93.900 133.200 94.000 ;
        RECT 131.000 93.600 133.200 93.900 ;
        RECT 131.000 93.500 131.400 93.600 ;
        RECT 134.200 93.200 134.600 94.600 ;
        RECT 137.100 94.300 139.000 94.700 ;
        RECT 137.100 93.700 137.500 94.300 ;
        RECT 139.300 94.000 139.600 95.000 ;
        RECT 131.000 93.100 131.400 93.200 ;
        RECT 126.100 92.700 127.400 93.100 ;
        RECT 129.100 92.800 131.400 93.100 ;
        RECT 134.100 92.800 134.600 93.200 ;
        RECT 136.600 93.400 137.500 93.700 ;
        RECT 139.000 93.700 139.600 94.000 ;
        RECT 136.600 93.100 137.000 93.400 ;
        RECT 127.000 91.100 127.400 92.700 ;
        RECT 135.800 92.700 137.000 93.100 ;
        RECT 127.800 91.100 128.200 92.500 ;
        RECT 128.600 91.100 129.000 92.500 ;
        RECT 129.400 91.100 129.800 92.500 ;
        RECT 131.000 91.100 131.400 92.500 ;
        RECT 132.600 91.100 133.000 92.500 ;
        RECT 133.400 91.100 133.800 92.500 ;
        RECT 134.200 91.100 134.600 92.500 ;
        RECT 135.000 91.100 135.400 92.500 ;
        RECT 135.800 91.100 136.200 92.700 ;
        RECT 139.000 91.100 139.400 93.700 ;
        RECT 139.900 93.400 140.300 95.600 ;
        RECT 142.200 95.600 142.500 95.900 ;
        RECT 142.200 95.200 142.800 95.600 ;
        RECT 140.600 95.100 141.000 95.200 ;
        RECT 141.400 95.100 141.800 95.200 ;
        RECT 140.600 94.800 141.800 95.100 ;
        RECT 141.400 94.400 141.800 94.800 ;
        RECT 142.200 93.700 142.500 95.200 ;
        RECT 144.700 94.200 145.000 95.900 ;
        RECT 147.000 95.600 147.300 95.900 ;
        RECT 145.400 94.800 145.800 95.600 ;
        RECT 147.000 95.200 147.600 95.600 ;
        RECT 146.200 94.400 146.600 95.200 ;
        RECT 144.600 93.800 145.000 94.200 ;
        RECT 139.800 93.000 140.300 93.400 ;
        RECT 141.400 93.400 142.500 93.700 ;
        RECT 139.800 91.100 140.200 93.000 ;
        RECT 141.400 91.100 141.800 93.400 ;
        RECT 143.800 92.400 144.200 93.200 ;
        RECT 144.700 92.100 145.000 93.800 ;
        RECT 147.000 93.700 147.300 95.200 ;
        RECT 144.600 91.100 145.000 92.100 ;
        RECT 146.200 93.400 147.300 93.700 ;
        RECT 146.200 91.100 146.600 93.400 ;
        RECT 148.600 92.400 149.000 93.200 ;
        RECT 149.400 91.100 149.800 99.900 ;
        RECT 2.200 87.900 2.600 89.900 ;
        RECT 2.900 88.200 3.300 88.600 ;
        RECT 1.400 86.400 1.800 87.200 ;
        RECT 0.600 86.100 1.000 86.200 ;
        RECT 2.200 86.100 2.500 87.900 ;
        RECT 3.000 87.800 3.400 88.200 ;
        RECT 3.800 87.900 4.200 89.900 ;
        RECT 4.600 88.000 5.000 89.900 ;
        RECT 6.200 88.000 6.600 89.900 ;
        RECT 4.600 87.900 6.600 88.000 ;
        RECT 7.600 89.200 8.000 89.900 ;
        RECT 7.600 88.800 8.200 89.200 ;
        RECT 3.900 87.200 4.200 87.900 ;
        RECT 4.700 87.700 6.500 87.900 ;
        RECT 5.800 87.200 6.200 87.400 ;
        RECT 3.800 86.800 5.100 87.200 ;
        RECT 5.800 86.900 6.600 87.200 ;
        RECT 7.600 87.100 8.000 88.800 ;
        RECT 10.300 88.200 10.700 88.600 ;
        RECT 10.200 87.800 10.600 88.200 ;
        RECT 11.000 87.900 11.400 89.900 ;
        RECT 6.200 86.800 6.600 86.900 ;
        RECT 7.100 86.900 8.000 87.100 ;
        RECT 7.100 86.800 7.900 86.900 ;
        RECT 3.000 86.100 3.400 86.200 ;
        RECT 0.600 85.800 1.400 86.100 ;
        RECT 2.200 85.800 3.400 86.100 ;
        RECT 1.000 85.600 1.400 85.800 ;
        RECT 3.000 85.100 3.300 85.800 ;
        RECT 3.800 85.100 4.200 85.200 ;
        RECT 4.800 85.100 5.100 86.800 ;
        RECT 5.400 85.800 5.800 86.600 ;
        RECT 7.100 85.200 7.400 86.800 ;
        RECT 8.200 85.800 9.000 86.200 ;
        RECT 10.200 86.100 10.600 86.200 ;
        RECT 11.100 86.100 11.400 87.900 ;
        RECT 14.000 89.200 14.400 89.900 ;
        RECT 14.000 88.800 14.600 89.200 ;
        RECT 11.800 86.400 12.200 87.200 ;
        RECT 14.000 87.100 14.400 88.800 ;
        RECT 18.400 87.200 18.800 89.900 ;
        RECT 19.800 87.900 20.200 89.900 ;
        RECT 22.000 88.100 22.800 89.900 ;
        RECT 19.800 87.600 21.100 87.900 ;
        RECT 20.700 87.500 21.100 87.600 ;
        RECT 21.400 87.400 22.200 87.800 ;
        RECT 13.500 86.900 14.400 87.100 ;
        RECT 18.200 87.100 18.800 87.200 ;
        RECT 19.800 87.100 20.600 87.200 ;
        RECT 22.500 87.100 22.800 88.100 ;
        RECT 24.600 87.900 25.000 89.900 ;
        RECT 25.700 89.200 26.100 89.900 ;
        RECT 25.400 88.800 26.100 89.200 ;
        RECT 25.700 88.200 26.100 88.800 ;
        RECT 25.700 87.900 26.600 88.200 ;
        RECT 27.800 87.900 28.200 89.900 ;
        RECT 28.600 88.000 29.000 89.900 ;
        RECT 30.200 88.000 30.600 89.900 ;
        RECT 28.600 87.900 30.600 88.000 ;
        RECT 31.000 87.900 31.400 89.900 ;
        RECT 31.800 88.000 32.200 89.900 ;
        RECT 33.400 88.000 33.800 89.900 ;
        RECT 31.800 87.900 33.800 88.000 ;
        RECT 23.100 87.400 23.500 87.800 ;
        RECT 23.800 87.600 25.000 87.900 ;
        RECT 23.800 87.500 24.200 87.600 ;
        RECT 13.500 86.800 14.300 86.900 ;
        RECT 18.200 86.800 19.300 87.100 ;
        RECT 19.800 87.000 20.900 87.100 ;
        RECT 19.800 86.800 22.000 87.000 ;
        RECT 12.600 86.100 13.000 86.200 ;
        RECT 10.200 85.800 11.400 86.100 ;
        RECT 12.200 85.800 13.000 86.100 ;
        RECT 0.600 84.800 2.600 85.100 ;
        RECT 0.600 81.100 1.000 84.800 ;
        RECT 2.200 81.100 2.600 84.800 ;
        RECT 3.000 81.100 3.400 85.100 ;
        RECT 3.800 84.800 4.500 85.100 ;
        RECT 4.800 84.800 5.300 85.100 ;
        RECT 7.000 84.800 7.400 85.200 ;
        RECT 9.400 84.800 9.800 85.600 ;
        RECT 10.300 85.100 10.600 85.800 ;
        RECT 12.200 85.600 12.600 85.800 ;
        RECT 13.500 85.200 13.800 86.800 ;
        RECT 14.600 85.800 15.400 86.200 ;
        RECT 17.400 85.800 18.200 86.200 ;
        RECT 4.200 84.200 4.500 84.800 ;
        RECT 4.200 83.800 4.600 84.200 ;
        RECT 4.900 81.100 5.300 84.800 ;
        RECT 7.100 83.500 7.400 84.800 ;
        RECT 7.800 83.800 8.200 84.600 ;
        RECT 7.100 83.200 8.900 83.500 ;
        RECT 7.100 83.100 7.400 83.200 ;
        RECT 7.000 81.100 7.400 83.100 ;
        RECT 8.600 83.100 8.900 83.200 ;
        RECT 8.600 81.100 9.000 83.100 ;
        RECT 10.200 81.100 10.600 85.100 ;
        RECT 11.000 84.800 13.000 85.100 ;
        RECT 13.400 84.800 13.800 85.200 ;
        RECT 15.800 84.800 16.200 85.600 ;
        RECT 16.600 84.800 17.000 85.600 ;
        RECT 19.000 85.200 19.300 86.800 ;
        RECT 20.600 86.700 22.000 86.800 ;
        RECT 21.600 86.600 22.000 86.700 ;
        RECT 22.300 86.800 22.800 87.100 ;
        RECT 23.200 87.200 23.500 87.400 ;
        RECT 23.200 86.800 23.600 87.200 ;
        RECT 24.200 86.800 25.000 87.200 ;
        RECT 22.300 86.200 22.600 86.800 ;
        RECT 20.900 86.100 21.300 86.200 ;
        RECT 20.900 85.800 21.700 86.100 ;
        RECT 22.200 85.800 22.600 86.200 ;
        RECT 21.300 85.700 21.700 85.800 ;
        RECT 19.000 84.800 19.400 85.200 ;
        RECT 22.300 85.100 22.600 85.800 ;
        RECT 25.400 85.800 25.800 86.200 ;
        RECT 25.400 85.200 25.700 85.800 ;
        RECT 19.800 84.800 21.100 85.100 ;
        RECT 11.000 81.100 11.400 84.800 ;
        RECT 12.600 81.100 13.000 84.800 ;
        RECT 13.500 83.500 13.800 84.800 ;
        RECT 14.200 84.100 14.600 84.600 ;
        RECT 15.800 84.100 16.200 84.200 ;
        RECT 14.200 83.800 16.200 84.100 ;
        RECT 18.200 83.800 18.600 84.600 ;
        RECT 19.000 83.500 19.300 84.800 ;
        RECT 13.500 83.200 15.300 83.500 ;
        RECT 13.500 83.100 13.800 83.200 ;
        RECT 13.400 81.100 13.800 83.100 ;
        RECT 15.000 83.100 15.300 83.200 ;
        RECT 17.500 83.200 19.300 83.500 ;
        RECT 17.500 83.100 17.800 83.200 ;
        RECT 15.000 81.100 15.400 83.100 ;
        RECT 17.400 81.100 17.800 83.100 ;
        RECT 19.000 83.100 19.300 83.200 ;
        RECT 19.000 81.100 19.400 83.100 ;
        RECT 19.800 81.100 20.200 84.800 ;
        RECT 20.700 84.700 21.100 84.800 ;
        RECT 22.000 81.100 22.800 85.100 ;
        RECT 23.800 84.800 25.000 85.100 ;
        RECT 23.800 84.700 24.200 84.800 ;
        RECT 24.600 81.100 25.000 84.800 ;
        RECT 25.400 84.400 25.800 85.200 ;
        RECT 26.200 81.100 26.600 87.900 ;
        RECT 27.000 86.800 27.400 87.600 ;
        RECT 27.900 87.200 28.200 87.900 ;
        RECT 28.700 87.700 30.500 87.900 ;
        RECT 29.800 87.200 30.200 87.400 ;
        RECT 31.100 87.200 31.400 87.900 ;
        RECT 31.900 87.700 33.700 87.900 ;
        RECT 33.000 87.200 33.400 87.400 ;
        RECT 27.800 86.800 29.100 87.200 ;
        RECT 29.800 86.900 30.600 87.200 ;
        RECT 30.200 86.800 30.600 86.900 ;
        RECT 31.000 86.800 32.300 87.200 ;
        RECT 33.000 86.900 33.800 87.200 ;
        RECT 34.800 87.100 35.200 89.900 ;
        RECT 37.500 88.200 37.900 88.600 ;
        RECT 37.400 87.800 37.800 88.200 ;
        RECT 38.200 87.900 38.600 89.900 ;
        RECT 40.900 88.200 41.300 89.900 ;
        RECT 43.300 89.200 43.700 89.900 ;
        RECT 43.300 88.800 44.200 89.200 ;
        RECT 43.300 88.200 43.700 88.800 ;
        RECT 33.400 86.800 33.800 86.900 ;
        RECT 34.300 86.900 35.200 87.100 ;
        RECT 37.400 87.100 37.800 87.200 ;
        RECT 38.300 87.100 38.600 87.900 ;
        RECT 40.600 87.800 41.800 88.200 ;
        RECT 43.300 87.900 44.200 88.200 ;
        RECT 45.400 87.900 45.800 89.900 ;
        RECT 46.200 88.000 46.600 89.900 ;
        RECT 47.800 88.000 48.200 89.900 ;
        RECT 51.500 89.200 51.900 89.900 ;
        RECT 51.000 88.800 51.900 89.200 ;
        RECT 51.500 88.200 51.900 88.800 ;
        RECT 46.200 87.900 48.200 88.000 ;
        RECT 51.000 87.900 51.900 88.200 ;
        RECT 52.600 88.000 53.000 89.900 ;
        RECT 54.200 88.000 54.600 89.900 ;
        RECT 52.600 87.900 54.600 88.000 ;
        RECT 55.000 87.900 55.400 89.900 ;
        RECT 57.400 87.900 57.800 89.900 ;
        RECT 59.300 89.200 59.700 89.900 ;
        RECT 59.000 88.800 59.700 89.200 ;
        RECT 58.100 88.200 58.500 88.600 ;
        RECT 59.300 88.200 59.700 88.800 ;
        RECT 61.700 88.200 62.100 89.900 ;
        RECT 40.600 87.200 40.900 87.800 ;
        RECT 34.300 86.800 35.100 86.900 ;
        RECT 37.400 86.800 38.600 87.100 ;
        RECT 27.000 86.200 27.300 86.800 ;
        RECT 28.800 86.200 29.100 86.800 ;
        RECT 27.000 85.800 27.400 86.200 ;
        RECT 28.600 85.800 29.100 86.200 ;
        RECT 29.400 86.100 29.800 86.600 ;
        RECT 30.200 86.100 30.600 86.200 ;
        RECT 29.400 85.800 30.600 86.100 ;
        RECT 27.800 85.100 28.200 85.200 ;
        RECT 28.800 85.100 29.100 85.800 ;
        RECT 31.000 85.100 31.400 85.200 ;
        RECT 32.000 85.100 32.300 86.800 ;
        RECT 32.600 85.800 33.000 86.600 ;
        RECT 34.300 85.200 34.600 86.800 ;
        RECT 35.400 85.800 36.200 86.200 ;
        RECT 37.400 86.100 37.800 86.200 ;
        RECT 38.300 86.100 38.600 86.800 ;
        RECT 39.000 86.400 39.400 87.200 ;
        RECT 40.600 86.800 41.000 87.200 ;
        RECT 39.800 86.100 40.200 86.200 ;
        RECT 37.400 85.800 38.600 86.100 ;
        RECT 39.400 85.800 40.200 86.100 ;
        RECT 27.800 84.800 28.500 85.100 ;
        RECT 28.800 84.800 29.300 85.100 ;
        RECT 31.000 84.800 31.700 85.100 ;
        RECT 32.000 84.800 32.500 85.100 ;
        RECT 34.200 84.800 34.600 85.200 ;
        RECT 36.600 84.800 37.000 85.600 ;
        RECT 37.500 85.100 37.800 85.800 ;
        RECT 39.400 85.600 39.800 85.800 ;
        RECT 28.200 84.200 28.500 84.800 ;
        RECT 28.200 83.800 28.600 84.200 ;
        RECT 28.900 81.100 29.300 84.800 ;
        RECT 31.400 84.200 31.700 84.800 ;
        RECT 32.100 84.200 32.500 84.800 ;
        RECT 31.400 83.800 31.800 84.200 ;
        RECT 32.100 83.800 33.000 84.200 ;
        RECT 32.100 81.100 32.500 83.800 ;
        RECT 34.300 83.500 34.600 84.800 ;
        RECT 35.000 83.800 35.400 84.600 ;
        RECT 34.300 83.200 36.100 83.500 ;
        RECT 34.300 83.100 34.600 83.200 ;
        RECT 34.200 81.100 34.600 83.100 ;
        RECT 35.800 83.100 36.100 83.200 ;
        RECT 35.800 81.100 36.200 83.100 ;
        RECT 37.400 81.100 37.800 85.100 ;
        RECT 38.200 84.800 40.200 85.100 ;
        RECT 38.200 81.100 38.600 84.800 ;
        RECT 39.800 81.100 40.200 84.800 ;
        RECT 41.400 81.100 41.800 87.800 ;
        RECT 43.000 84.400 43.400 85.200 ;
        RECT 43.800 81.100 44.200 87.900 ;
        RECT 44.600 86.800 45.000 87.600 ;
        RECT 45.500 87.200 45.800 87.900 ;
        RECT 46.300 87.700 48.100 87.900 ;
        RECT 47.400 87.200 47.800 87.400 ;
        RECT 45.400 86.800 46.700 87.200 ;
        RECT 47.400 86.900 48.200 87.200 ;
        RECT 47.800 86.800 48.200 86.900 ;
        RECT 50.200 86.800 50.600 87.600 ;
        RECT 44.600 86.100 45.000 86.200 ;
        RECT 46.400 86.100 46.700 86.800 ;
        RECT 44.600 85.800 46.700 86.100 ;
        RECT 47.000 86.100 47.400 86.600 ;
        RECT 47.800 86.100 48.200 86.200 ;
        RECT 47.000 85.800 48.200 86.100 ;
        RECT 45.400 85.100 45.800 85.200 ;
        RECT 46.400 85.100 46.700 85.800 ;
        RECT 45.400 84.800 46.100 85.100 ;
        RECT 46.400 84.800 46.900 85.100 ;
        RECT 45.800 84.200 46.100 84.800 ;
        RECT 45.800 83.800 46.200 84.200 ;
        RECT 46.500 81.100 46.900 84.800 ;
        RECT 51.000 81.100 51.400 87.900 ;
        RECT 52.700 87.700 54.500 87.900 ;
        RECT 53.000 87.200 53.400 87.400 ;
        RECT 55.000 87.200 55.300 87.900 ;
        RECT 57.400 87.200 57.700 87.900 ;
        RECT 58.200 87.800 58.600 88.200 ;
        RECT 59.300 87.900 60.200 88.200 ;
        RECT 52.600 86.900 53.400 87.200 ;
        RECT 52.600 86.800 53.000 86.900 ;
        RECT 54.100 86.800 55.400 87.200 ;
        RECT 57.400 86.800 57.800 87.200 ;
        RECT 52.600 86.100 53.000 86.200 ;
        RECT 53.400 86.100 53.800 86.600 ;
        RECT 52.600 85.800 53.800 86.100 ;
        RECT 51.800 84.400 52.200 85.200 ;
        RECT 54.100 85.100 54.400 86.800 ;
        RECT 57.400 86.100 57.700 86.800 ;
        RECT 58.200 86.100 58.600 86.200 ;
        RECT 57.400 85.800 58.600 86.100 ;
        RECT 55.000 85.100 55.400 85.200 ;
        RECT 58.200 85.100 58.500 85.800 ;
        RECT 53.900 84.800 54.400 85.100 ;
        RECT 54.700 84.800 55.400 85.100 ;
        RECT 55.800 84.800 57.800 85.100 ;
        RECT 53.900 84.200 54.300 84.800 ;
        RECT 54.700 84.200 55.000 84.800 ;
        RECT 53.400 83.800 54.300 84.200 ;
        RECT 54.600 83.800 55.000 84.200 ;
        RECT 53.900 81.100 54.300 83.800 ;
        RECT 55.800 81.100 56.200 84.800 ;
        RECT 57.400 81.100 57.800 84.800 ;
        RECT 58.200 81.100 58.600 85.100 ;
        RECT 59.800 81.100 60.200 87.900 ;
        RECT 61.400 87.800 62.600 88.200 ;
        RECT 63.800 87.900 64.200 89.900 ;
        RECT 64.600 88.000 65.000 89.900 ;
        RECT 66.200 88.000 66.600 89.900 ;
        RECT 64.600 87.900 66.600 88.000 ;
        RECT 67.000 87.900 67.400 89.900 ;
        RECT 67.800 88.000 68.200 89.900 ;
        RECT 69.400 88.000 69.800 89.900 ;
        RECT 67.800 87.900 69.800 88.000 ;
        RECT 70.200 88.000 70.600 89.900 ;
        RECT 71.800 88.000 72.200 89.900 ;
        RECT 70.200 87.900 72.200 88.000 ;
        RECT 72.600 87.900 73.000 89.900 ;
        RECT 73.700 89.200 74.100 89.900 ;
        RECT 73.400 88.800 74.100 89.200 ;
        RECT 73.700 88.200 74.100 88.800 ;
        RECT 73.700 87.900 74.600 88.200 ;
        RECT 61.400 87.200 61.700 87.800 ;
        RECT 61.400 86.800 61.800 87.200 ;
        RECT 62.200 81.100 62.600 87.800 ;
        RECT 63.900 87.200 64.200 87.900 ;
        RECT 64.700 87.700 66.500 87.900 ;
        RECT 65.800 87.200 66.200 87.400 ;
        RECT 67.100 87.200 67.400 87.900 ;
        RECT 67.900 87.700 69.700 87.900 ;
        RECT 70.300 87.700 72.100 87.900 ;
        RECT 69.000 87.200 69.400 87.400 ;
        RECT 70.600 87.200 71.000 87.400 ;
        RECT 72.600 87.200 72.900 87.900 ;
        RECT 63.800 86.800 65.100 87.200 ;
        RECT 65.800 86.900 66.600 87.200 ;
        RECT 66.200 86.800 66.600 86.900 ;
        RECT 67.000 86.800 68.300 87.200 ;
        RECT 69.000 87.100 69.800 87.200 ;
        RECT 70.200 87.100 71.000 87.200 ;
        RECT 69.000 86.900 71.000 87.100 ;
        RECT 69.400 86.800 70.600 86.900 ;
        RECT 71.700 86.800 73.000 87.200 ;
        RECT 63.800 85.100 64.200 85.200 ;
        RECT 64.800 85.100 65.100 86.800 ;
        RECT 65.400 85.800 65.800 86.600 ;
        RECT 67.000 85.100 67.400 85.200 ;
        RECT 68.000 85.100 68.300 86.800 ;
        RECT 68.600 86.100 69.000 86.600 ;
        RECT 69.400 86.100 69.800 86.200 ;
        RECT 71.000 86.100 71.400 86.600 ;
        RECT 68.600 85.800 71.400 86.100 ;
        RECT 71.700 85.100 72.000 86.800 ;
        RECT 72.600 85.100 73.000 85.200 ;
        RECT 63.800 84.800 64.500 85.100 ;
        RECT 64.800 84.800 65.300 85.100 ;
        RECT 67.000 84.800 67.700 85.100 ;
        RECT 68.000 84.800 68.500 85.100 ;
        RECT 64.200 84.200 64.500 84.800 ;
        RECT 64.200 83.800 64.600 84.200 ;
        RECT 64.900 81.100 65.300 84.800 ;
        RECT 67.400 84.200 67.700 84.800 ;
        RECT 67.400 83.800 67.800 84.200 ;
        RECT 68.100 81.100 68.500 84.800 ;
        RECT 71.500 84.800 72.000 85.100 ;
        RECT 72.300 84.800 73.000 85.100 ;
        RECT 71.500 81.100 71.900 84.800 ;
        RECT 72.300 84.200 72.600 84.800 ;
        RECT 72.200 83.800 72.600 84.200 ;
        RECT 74.200 81.100 74.600 87.900 ;
        RECT 75.800 87.900 76.200 89.900 ;
        RECT 78.000 89.200 78.800 89.900 ;
        RECT 78.000 88.800 79.400 89.200 ;
        RECT 78.000 88.100 78.800 88.800 ;
        RECT 75.800 87.600 77.000 87.900 ;
        RECT 76.600 87.500 77.000 87.600 ;
        RECT 77.300 87.400 77.700 87.800 ;
        RECT 77.300 87.200 77.600 87.400 ;
        RECT 75.800 86.800 76.600 87.200 ;
        RECT 77.200 86.800 77.600 87.200 ;
        RECT 78.000 87.100 78.300 88.100 ;
        RECT 80.600 87.900 81.000 89.900 ;
        RECT 81.400 87.900 81.800 89.900 ;
        RECT 83.500 89.200 83.900 89.900 ;
        RECT 83.500 88.800 84.200 89.200 ;
        RECT 83.500 88.400 83.900 88.800 ;
        RECT 83.500 87.900 84.200 88.400 ;
        RECT 78.600 87.400 79.400 87.800 ;
        RECT 79.700 87.600 81.000 87.900 ;
        RECT 81.500 87.800 81.800 87.900 ;
        RECT 81.500 87.600 82.400 87.800 ;
        RECT 79.700 87.500 80.100 87.600 ;
        RECT 81.500 87.500 83.600 87.600 ;
        RECT 82.100 87.300 83.600 87.500 ;
        RECT 83.200 87.200 83.600 87.300 ;
        RECT 80.200 87.100 81.000 87.200 ;
        RECT 81.400 87.100 81.800 87.200 ;
        RECT 78.000 86.800 78.500 87.100 ;
        RECT 79.900 87.000 81.800 87.100 ;
        RECT 78.200 86.200 78.500 86.800 ;
        RECT 78.800 86.800 81.800 87.000 ;
        RECT 82.400 86.900 82.800 87.000 ;
        RECT 78.800 86.700 80.200 86.800 ;
        RECT 78.800 86.600 79.200 86.700 ;
        RECT 81.400 86.400 81.800 86.800 ;
        RECT 82.300 86.600 82.800 86.900 ;
        RECT 82.300 86.200 82.600 86.600 ;
        RECT 78.200 85.800 78.600 86.200 ;
        RECT 79.500 86.100 79.900 86.200 ;
        RECT 79.100 85.800 79.900 86.100 ;
        RECT 82.200 85.800 82.600 86.200 ;
        RECT 78.200 85.100 78.500 85.800 ;
        RECT 79.100 85.700 79.500 85.800 ;
        RECT 83.200 85.500 83.500 87.200 ;
        RECT 83.900 86.200 84.200 87.900 ;
        RECT 83.800 85.800 84.200 86.200 ;
        RECT 82.300 85.200 83.500 85.500 ;
        RECT 75.800 84.800 77.000 85.100 ;
        RECT 75.800 81.100 76.200 84.800 ;
        RECT 76.600 84.700 77.000 84.800 ;
        RECT 78.000 81.100 78.800 85.100 ;
        RECT 79.700 84.800 81.000 85.100 ;
        RECT 79.700 84.700 80.100 84.800 ;
        RECT 80.600 81.100 81.000 84.800 ;
        RECT 82.300 83.100 82.600 85.200 ;
        RECT 83.900 85.100 84.200 85.800 ;
        RECT 82.200 81.100 82.600 83.100 ;
        RECT 83.800 81.100 84.200 85.100 ;
        RECT 84.600 81.100 85.000 89.900 ;
        RECT 87.000 81.100 87.400 89.900 ;
        RECT 88.600 88.000 89.000 89.900 ;
        RECT 90.200 88.000 90.600 89.900 ;
        RECT 88.600 87.900 90.600 88.000 ;
        RECT 91.000 87.900 91.400 89.900 ;
        RECT 91.900 88.200 92.300 88.600 ;
        RECT 88.700 87.700 90.500 87.900 ;
        RECT 89.000 87.200 89.400 87.400 ;
        RECT 91.000 87.200 91.300 87.900 ;
        RECT 91.800 87.800 92.200 88.200 ;
        RECT 92.600 87.900 93.000 89.900 ;
        RECT 95.800 88.900 96.200 89.900 ;
        RECT 88.600 86.900 89.400 87.200 ;
        RECT 90.100 87.100 91.400 87.200 ;
        RECT 91.800 87.100 92.200 87.200 ;
        RECT 88.600 86.800 89.000 86.900 ;
        RECT 90.100 86.800 92.200 87.100 ;
        RECT 89.400 85.800 89.800 86.600 ;
        RECT 90.100 85.100 90.400 86.800 ;
        RECT 91.800 86.100 92.200 86.200 ;
        RECT 92.700 86.100 93.000 87.900 ;
        RECT 95.000 87.800 95.400 88.600 ;
        RECT 95.900 88.100 96.200 88.900 ;
        RECT 97.400 88.100 97.800 88.600 ;
        RECT 95.800 87.800 97.800 88.100 ;
        RECT 95.900 87.200 96.200 87.800 ;
        RECT 93.400 86.400 93.800 87.200 ;
        RECT 95.800 86.800 96.200 87.200 ;
        RECT 94.200 86.100 94.600 86.200 ;
        RECT 95.900 86.100 96.200 86.800 ;
        RECT 98.200 87.100 98.600 89.900 ;
        RECT 100.600 87.900 101.000 89.900 ;
        RECT 102.800 89.200 103.600 89.900 ;
        RECT 102.200 88.800 103.600 89.200 ;
        RECT 102.800 88.100 103.600 88.800 ;
        RECT 100.600 87.600 101.800 87.900 ;
        RECT 101.400 87.500 101.800 87.600 ;
        RECT 102.100 87.400 102.500 87.800 ;
        RECT 102.100 87.200 102.400 87.400 ;
        RECT 100.600 87.100 101.400 87.200 ;
        RECT 98.200 86.800 101.400 87.100 ;
        RECT 102.000 86.800 102.400 87.200 ;
        RECT 91.800 85.800 93.000 86.100 ;
        RECT 93.800 85.800 96.200 86.100 ;
        RECT 91.000 85.100 91.400 85.200 ;
        RECT 91.900 85.100 92.200 85.800 ;
        RECT 93.800 85.600 94.200 85.800 ;
        RECT 95.900 85.100 96.200 85.800 ;
        RECT 96.600 85.400 97.000 86.200 ;
        RECT 89.900 84.800 90.400 85.100 ;
        RECT 90.700 84.800 91.400 85.100 ;
        RECT 89.900 81.100 90.300 84.800 ;
        RECT 90.700 84.200 91.000 84.800 ;
        RECT 90.600 83.800 91.000 84.200 ;
        RECT 91.800 81.100 92.200 85.100 ;
        RECT 92.600 84.800 94.600 85.100 ;
        RECT 92.600 81.100 93.000 84.800 ;
        RECT 94.200 81.100 94.600 84.800 ;
        RECT 95.800 84.700 96.700 85.100 ;
        RECT 96.300 81.100 96.700 84.700 ;
        RECT 98.200 81.100 98.600 86.800 ;
        RECT 102.800 86.400 103.100 88.100 ;
        RECT 105.400 87.900 105.800 89.900 ;
        RECT 106.500 89.200 106.900 89.900 ;
        RECT 106.200 88.800 106.900 89.200 ;
        RECT 106.500 88.200 106.900 88.800 ;
        RECT 106.500 87.900 107.400 88.200 ;
        RECT 103.400 87.700 104.200 87.800 ;
        RECT 103.400 87.400 104.400 87.700 ;
        RECT 104.700 87.600 105.800 87.900 ;
        RECT 104.700 87.500 105.100 87.600 ;
        RECT 104.100 87.200 104.400 87.400 ;
        RECT 103.400 86.700 103.800 87.100 ;
        RECT 104.100 86.900 105.800 87.200 ;
        RECT 105.000 86.800 105.800 86.900 ;
        RECT 102.600 86.200 103.100 86.400 ;
        RECT 102.200 86.100 103.100 86.200 ;
        RECT 103.500 86.400 103.800 86.700 ;
        RECT 103.500 86.100 104.800 86.400 ;
        RECT 102.200 85.800 102.900 86.100 ;
        RECT 104.400 86.000 104.800 86.100 ;
        RECT 102.600 85.100 102.900 85.800 ;
        RECT 103.300 85.700 103.700 85.800 ;
        RECT 103.300 85.400 105.000 85.700 ;
        RECT 104.700 85.100 105.000 85.400 ;
        RECT 100.600 84.800 101.800 85.100 ;
        RECT 102.600 84.800 103.600 85.100 ;
        RECT 100.600 81.100 101.000 84.800 ;
        RECT 101.400 84.700 101.800 84.800 ;
        RECT 102.800 81.100 103.600 84.800 ;
        RECT 104.700 84.800 105.800 85.100 ;
        RECT 104.700 84.700 105.100 84.800 ;
        RECT 105.400 81.100 105.800 84.800 ;
        RECT 107.000 81.100 107.400 87.900 ;
        RECT 107.800 86.800 108.200 87.600 ;
        RECT 109.400 81.100 109.800 89.900 ;
        RECT 112.600 87.900 113.000 89.900 ;
        RECT 113.300 88.200 113.700 88.600 ;
        RECT 113.400 88.100 113.800 88.200 ;
        RECT 114.200 88.100 114.600 89.900 ;
        RECT 110.200 86.800 110.600 87.600 ;
        RECT 111.800 86.400 112.200 87.200 ;
        RECT 111.000 86.100 111.400 86.200 ;
        RECT 112.600 86.100 112.900 87.900 ;
        RECT 113.400 87.800 114.600 88.100 ;
        RECT 115.000 88.000 115.400 89.900 ;
        RECT 116.600 88.000 117.000 89.900 ;
        RECT 118.200 88.900 118.600 89.900 ;
        RECT 120.600 88.900 121.000 89.900 ;
        RECT 115.000 87.900 117.000 88.000 ;
        RECT 117.400 88.100 117.800 88.200 ;
        RECT 118.200 88.100 118.500 88.900 ;
        RECT 114.300 87.200 114.600 87.800 ;
        RECT 115.100 87.700 116.900 87.900 ;
        RECT 117.400 87.800 118.500 88.100 ;
        RECT 119.000 87.800 119.400 88.600 ;
        RECT 119.800 87.800 120.200 88.600 ;
        RECT 120.700 87.800 121.000 88.900 ;
        RECT 122.200 87.900 122.600 89.900 ;
        RECT 116.200 87.200 116.600 87.400 ;
        RECT 118.200 87.200 118.500 87.800 ;
        RECT 120.700 87.500 121.900 87.800 ;
        RECT 114.200 86.800 115.500 87.200 ;
        RECT 116.200 87.100 117.000 87.200 ;
        RECT 116.200 86.900 117.700 87.100 ;
        RECT 116.600 86.800 117.700 86.900 ;
        RECT 113.400 86.100 113.800 86.200 ;
        RECT 111.000 85.800 111.800 86.100 ;
        RECT 112.600 85.800 113.800 86.100 ;
        RECT 111.400 85.600 111.800 85.800 ;
        RECT 113.400 85.100 113.700 85.800 ;
        RECT 114.200 85.100 114.600 85.200 ;
        RECT 115.200 85.100 115.500 86.800 ;
        RECT 115.800 86.100 116.200 86.600 ;
        RECT 117.400 86.200 117.700 86.800 ;
        RECT 118.200 86.800 118.600 87.200 ;
        RECT 120.600 86.800 121.100 87.200 ;
        RECT 116.600 86.100 117.000 86.200 ;
        RECT 115.800 85.800 117.000 86.100 ;
        RECT 117.400 85.400 117.800 86.200 ;
        RECT 118.200 85.100 118.500 86.800 ;
        RECT 120.800 86.400 121.200 86.800 ;
        RECT 121.600 86.000 121.900 87.500 ;
        RECT 122.300 87.100 122.600 87.900 ;
        RECT 124.600 87.900 125.000 89.900 ;
        RECT 125.300 88.200 125.700 88.600 ;
        RECT 123.000 87.100 123.400 87.200 ;
        RECT 122.200 86.800 123.400 87.100 ;
        RECT 122.300 86.200 122.600 86.800 ;
        RECT 123.800 86.400 124.200 87.200 ;
        RECT 121.500 85.700 121.900 86.000 ;
        RECT 122.200 85.800 122.600 86.200 ;
        RECT 123.000 86.100 123.400 86.200 ;
        RECT 124.600 86.100 124.900 87.900 ;
        RECT 125.400 87.800 125.800 88.200 ;
        RECT 126.200 88.000 126.600 89.900 ;
        RECT 127.800 88.000 128.200 89.900 ;
        RECT 126.200 87.900 128.200 88.000 ;
        RECT 128.600 87.900 129.000 89.900 ;
        RECT 129.400 88.000 129.800 89.900 ;
        RECT 131.000 88.000 131.400 89.900 ;
        RECT 129.400 87.900 131.400 88.000 ;
        RECT 131.800 87.900 132.200 89.900 ;
        RECT 132.600 87.900 133.000 89.900 ;
        RECT 134.800 88.100 135.600 89.900 ;
        RECT 126.300 87.700 128.100 87.900 ;
        RECT 126.600 87.200 127.000 87.400 ;
        RECT 128.600 87.200 128.900 87.900 ;
        RECT 129.500 87.700 131.300 87.900 ;
        RECT 129.800 87.200 130.200 87.400 ;
        RECT 131.800 87.200 132.100 87.900 ;
        RECT 132.600 87.600 133.700 87.900 ;
        RECT 134.200 87.700 135.000 87.800 ;
        RECT 133.300 87.500 133.700 87.600 ;
        RECT 134.000 87.400 135.000 87.700 ;
        RECT 134.000 87.200 134.300 87.400 ;
        RECT 126.200 86.900 127.000 87.200 ;
        RECT 126.200 86.800 126.600 86.900 ;
        RECT 127.700 86.800 129.000 87.200 ;
        RECT 129.400 86.900 130.200 87.200 ;
        RECT 129.400 86.800 129.800 86.900 ;
        RECT 130.900 86.800 132.200 87.200 ;
        RECT 132.600 86.900 134.300 87.200 ;
        RECT 132.600 86.800 133.400 86.900 ;
        RECT 125.400 86.100 125.800 86.200 ;
        RECT 123.000 85.800 123.800 86.100 ;
        RECT 124.600 85.800 125.800 86.100 ;
        RECT 127.000 85.800 127.400 86.600 ;
        RECT 119.800 85.600 121.900 85.700 ;
        RECT 119.800 85.400 121.800 85.600 ;
        RECT 111.000 84.800 113.000 85.100 ;
        RECT 111.000 81.100 111.400 84.800 ;
        RECT 112.600 81.100 113.000 84.800 ;
        RECT 113.400 81.100 113.800 85.100 ;
        RECT 114.200 84.800 114.900 85.100 ;
        RECT 115.200 84.800 115.700 85.100 ;
        RECT 114.600 84.200 114.900 84.800 ;
        RECT 114.600 83.800 115.000 84.200 ;
        RECT 115.300 81.100 115.700 84.800 ;
        RECT 117.700 84.700 118.600 85.100 ;
        RECT 117.700 81.100 118.100 84.700 ;
        RECT 119.800 81.100 120.200 85.400 ;
        RECT 122.300 85.100 122.600 85.800 ;
        RECT 123.400 85.600 123.800 85.800 ;
        RECT 125.400 85.100 125.700 85.800 ;
        RECT 127.700 85.100 128.000 86.800 ;
        RECT 128.600 86.100 129.000 86.200 ;
        RECT 130.200 86.100 130.600 86.600 ;
        RECT 128.600 85.800 130.600 86.100 ;
        RECT 128.600 85.100 129.000 85.200 ;
        RECT 130.900 85.100 131.200 86.800 ;
        RECT 134.600 86.700 135.000 87.100 ;
        RECT 134.600 86.400 134.900 86.700 ;
        RECT 133.600 86.100 134.900 86.400 ;
        RECT 135.300 86.400 135.600 88.100 ;
        RECT 137.400 87.900 137.800 89.900 ;
        RECT 135.900 87.400 136.300 87.800 ;
        RECT 136.600 87.600 137.800 87.900 ;
        RECT 139.800 87.900 140.200 89.900 ;
        RECT 140.500 88.200 140.900 88.600 ;
        RECT 136.600 87.500 137.000 87.600 ;
        RECT 136.000 87.200 136.300 87.400 ;
        RECT 136.000 86.800 136.400 87.200 ;
        RECT 137.000 86.800 137.800 87.200 ;
        RECT 139.000 86.400 139.400 87.200 ;
        RECT 135.300 86.200 135.800 86.400 ;
        RECT 135.300 86.100 136.200 86.200 ;
        RECT 133.600 86.000 134.000 86.100 ;
        RECT 135.500 85.800 136.200 86.100 ;
        RECT 138.200 86.100 138.600 86.200 ;
        RECT 139.800 86.100 140.100 87.900 ;
        RECT 140.600 87.800 141.000 88.200 ;
        RECT 141.400 87.900 141.800 89.900 ;
        RECT 142.200 88.000 142.600 89.900 ;
        RECT 143.800 88.000 144.200 89.900 ;
        RECT 142.200 87.900 144.200 88.000 ;
        RECT 141.500 87.200 141.800 87.900 ;
        RECT 142.300 87.700 144.100 87.900 ;
        RECT 143.400 87.200 143.800 87.400 ;
        RECT 141.400 86.800 142.700 87.200 ;
        RECT 143.400 87.100 144.200 87.200 ;
        RECT 144.600 87.100 145.000 89.900 ;
        RECT 145.400 87.800 145.800 88.600 ;
        RECT 146.200 87.600 146.600 89.900 ;
        RECT 148.900 88.200 149.300 89.900 ;
        RECT 148.900 87.900 149.800 88.200 ;
        RECT 146.200 87.300 147.300 87.600 ;
        RECT 143.400 86.900 145.000 87.100 ;
        RECT 143.800 86.800 145.000 86.900 ;
        RECT 140.600 86.100 141.000 86.200 ;
        RECT 138.200 85.800 139.000 86.100 ;
        RECT 139.800 85.800 141.000 86.100 ;
        RECT 134.700 85.700 135.100 85.800 ;
        RECT 133.400 85.400 135.100 85.700 ;
        RECT 131.800 85.100 132.200 85.200 ;
        RECT 133.400 85.100 133.700 85.400 ;
        RECT 135.500 85.100 135.800 85.800 ;
        RECT 138.600 85.600 139.000 85.800 ;
        RECT 140.600 85.100 140.900 85.800 ;
        RECT 141.400 85.100 141.800 85.200 ;
        RECT 142.400 85.100 142.700 86.800 ;
        RECT 121.900 84.800 122.600 85.100 ;
        RECT 123.000 84.800 125.000 85.100 ;
        RECT 121.900 81.100 122.300 84.800 ;
        RECT 123.000 81.100 123.400 84.800 ;
        RECT 124.600 81.100 125.000 84.800 ;
        RECT 125.400 81.100 125.800 85.100 ;
        RECT 127.500 84.800 128.000 85.100 ;
        RECT 128.300 84.800 129.000 85.100 ;
        RECT 130.700 84.800 131.200 85.100 ;
        RECT 131.500 84.800 132.200 85.100 ;
        RECT 132.600 84.800 133.700 85.100 ;
        RECT 127.500 81.100 127.900 84.800 ;
        RECT 128.300 84.200 128.600 84.800 ;
        RECT 128.200 83.800 128.600 84.200 ;
        RECT 130.700 81.100 131.100 84.800 ;
        RECT 131.500 84.200 131.800 84.800 ;
        RECT 131.400 83.800 131.800 84.200 ;
        RECT 132.600 81.100 133.000 84.800 ;
        RECT 133.300 84.700 133.700 84.800 ;
        RECT 134.800 84.800 135.800 85.100 ;
        RECT 136.600 84.800 137.800 85.100 ;
        RECT 134.800 81.100 135.600 84.800 ;
        RECT 136.600 84.700 137.000 84.800 ;
        RECT 137.400 81.100 137.800 84.800 ;
        RECT 138.200 84.800 140.200 85.100 ;
        RECT 138.200 81.100 138.600 84.800 ;
        RECT 139.800 81.100 140.200 84.800 ;
        RECT 140.600 81.100 141.000 85.100 ;
        RECT 141.400 84.800 142.100 85.100 ;
        RECT 142.400 84.800 142.900 85.100 ;
        RECT 141.800 84.200 142.100 84.800 ;
        RECT 141.800 83.800 142.200 84.200 ;
        RECT 142.500 81.100 142.900 84.800 ;
        RECT 144.600 81.100 145.000 86.800 ;
        RECT 146.200 85.800 146.600 86.600 ;
        RECT 147.000 85.800 147.300 87.300 ;
        RECT 147.000 85.400 147.600 85.800 ;
        RECT 147.000 85.100 147.300 85.400 ;
        RECT 146.200 84.800 147.300 85.100 ;
        RECT 146.200 81.100 146.600 84.800 ;
        RECT 148.600 84.400 149.000 85.200 ;
        RECT 149.400 81.100 149.800 87.900 ;
        RECT 150.200 86.800 150.600 87.600 ;
        RECT 0.600 77.900 1.000 79.900 ;
        RECT 0.700 77.800 1.000 77.900 ;
        RECT 2.200 77.900 2.600 79.900 ;
        RECT 2.200 77.800 2.500 77.900 ;
        RECT 0.700 77.500 2.500 77.800 ;
        RECT 0.700 76.200 1.000 77.500 ;
        RECT 1.400 76.400 1.800 77.200 ;
        RECT 4.200 76.800 4.600 77.200 ;
        RECT 4.200 76.200 4.500 76.800 ;
        RECT 4.900 76.200 5.300 79.900 ;
        RECT 7.000 77.900 7.400 79.900 ;
        RECT 7.100 77.800 7.400 77.900 ;
        RECT 8.600 77.900 9.000 79.900 ;
        RECT 8.600 77.800 8.900 77.900 ;
        RECT 7.100 77.500 8.900 77.800 ;
        RECT 7.100 76.200 7.400 77.500 ;
        RECT 7.800 76.400 8.200 77.200 ;
        RECT 0.600 75.800 1.000 76.200 ;
        RECT 0.700 74.200 1.000 75.800 ;
        RECT 3.000 75.400 3.400 76.200 ;
        RECT 3.800 75.900 4.500 76.200 ;
        RECT 4.800 75.900 5.300 76.200 ;
        RECT 3.800 75.800 4.200 75.900 ;
        RECT 3.800 75.200 4.100 75.800 ;
        RECT 1.800 74.800 2.600 75.200 ;
        RECT 3.800 74.800 4.200 75.200 ;
        RECT 4.800 74.200 5.100 75.900 ;
        RECT 7.000 75.800 7.400 76.200 ;
        RECT 5.400 74.400 5.800 75.200 ;
        RECT 7.100 74.200 7.400 75.800 ;
        RECT 9.400 75.400 9.800 76.200 ;
        RECT 10.200 75.900 10.600 79.900 ;
        RECT 11.000 76.200 11.400 79.900 ;
        RECT 12.600 76.200 13.000 79.900 ;
        RECT 14.200 77.900 14.600 79.900 ;
        RECT 14.300 77.800 14.600 77.900 ;
        RECT 15.800 77.900 16.200 79.900 ;
        RECT 15.800 77.800 16.100 77.900 ;
        RECT 14.300 77.500 16.100 77.800 ;
        RECT 15.000 76.400 15.400 77.200 ;
        RECT 15.800 76.200 16.100 77.500 ;
        RECT 11.000 75.900 13.000 76.200 ;
        RECT 10.300 75.200 10.600 75.900 ;
        RECT 13.400 75.400 13.800 76.200 ;
        RECT 15.800 75.800 16.200 76.200 ;
        RECT 16.600 75.800 17.000 76.600 ;
        RECT 12.200 75.200 12.600 75.400 ;
        RECT 8.200 74.800 9.000 75.200 ;
        RECT 10.200 74.900 11.400 75.200 ;
        RECT 12.200 74.900 13.000 75.200 ;
        RECT 10.200 74.800 10.600 74.900 ;
        RECT 0.700 74.100 1.500 74.200 ;
        RECT 0.700 73.900 1.600 74.100 ;
        RECT 1.200 71.100 1.600 73.900 ;
        RECT 3.800 73.800 5.100 74.200 ;
        RECT 6.200 74.100 6.600 74.200 ;
        RECT 5.800 73.800 6.600 74.100 ;
        RECT 7.100 74.100 7.900 74.200 ;
        RECT 7.100 73.900 8.000 74.100 ;
        RECT 3.900 73.100 4.200 73.800 ;
        RECT 5.800 73.600 6.200 73.800 ;
        RECT 4.700 73.100 6.500 73.300 ;
        RECT 3.800 71.100 4.200 73.100 ;
        RECT 4.600 73.000 6.600 73.100 ;
        RECT 4.600 71.100 5.000 73.000 ;
        RECT 6.200 71.100 6.600 73.000 ;
        RECT 7.600 71.100 8.000 73.900 ;
        RECT 10.200 72.800 10.600 73.200 ;
        RECT 11.100 73.100 11.400 74.900 ;
        RECT 12.600 74.800 13.000 74.900 ;
        RECT 14.200 74.800 15.000 75.200 ;
        RECT 11.800 73.800 12.200 74.600 ;
        RECT 15.800 74.200 16.100 75.800 ;
        RECT 15.300 74.100 16.100 74.200 ;
        RECT 15.200 73.900 16.100 74.100 ;
        RECT 10.300 72.400 10.700 72.800 ;
        RECT 11.000 71.100 11.400 73.100 ;
        RECT 15.200 71.100 15.600 73.900 ;
        RECT 17.400 73.100 17.800 79.900 ;
        RECT 20.300 76.200 20.700 79.900 ;
        RECT 21.000 76.800 21.400 77.200 ;
        RECT 21.100 76.200 21.400 76.800 ;
        RECT 23.500 76.200 23.900 79.900 ;
        RECT 24.200 76.800 24.600 77.200 ;
        RECT 24.300 76.200 24.600 76.800 ;
        RECT 19.800 75.800 20.800 76.200 ;
        RECT 21.100 75.900 21.800 76.200 ;
        RECT 23.500 75.900 24.000 76.200 ;
        RECT 24.300 75.900 25.000 76.200 ;
        RECT 21.400 75.800 21.800 75.900 ;
        RECT 19.800 74.400 20.200 75.200 ;
        RECT 20.500 74.200 20.800 75.800 ;
        RECT 23.000 74.400 23.400 75.200 ;
        RECT 23.700 75.100 24.000 75.900 ;
        RECT 24.600 75.800 25.000 75.900 ;
        RECT 25.400 75.800 25.800 76.600 ;
        RECT 25.400 75.100 25.700 75.800 ;
        RECT 23.700 74.800 25.700 75.100 ;
        RECT 23.700 74.200 24.000 74.800 ;
        RECT 18.200 73.400 18.600 74.200 ;
        RECT 19.000 74.100 19.400 74.200 ;
        RECT 19.000 73.800 19.800 74.100 ;
        RECT 20.500 73.800 21.800 74.200 ;
        RECT 22.200 74.100 22.600 74.200 ;
        RECT 22.200 73.800 23.000 74.100 ;
        RECT 23.700 73.800 25.000 74.200 ;
        RECT 19.400 73.600 19.800 73.800 ;
        RECT 19.100 73.100 20.900 73.300 ;
        RECT 21.400 73.100 21.700 73.800 ;
        RECT 22.600 73.600 23.000 73.800 ;
        RECT 22.300 73.100 24.100 73.300 ;
        RECT 24.600 73.100 24.900 73.800 ;
        RECT 26.200 73.100 26.600 79.900 ;
        RECT 27.800 76.100 28.200 76.200 ;
        RECT 28.600 76.100 29.000 79.900 ;
        RECT 29.800 76.800 30.200 77.200 ;
        RECT 29.800 76.200 30.100 76.800 ;
        RECT 30.500 76.200 30.900 79.900 ;
        RECT 33.900 76.200 34.300 79.900 ;
        RECT 34.600 76.800 35.000 77.200 ;
        RECT 34.700 76.200 35.000 76.800 ;
        RECT 29.400 76.100 30.100 76.200 ;
        RECT 27.800 75.900 30.100 76.100 ;
        RECT 30.400 75.900 30.900 76.200 ;
        RECT 27.800 75.800 29.800 75.900 ;
        RECT 27.000 73.400 27.400 74.200 ;
        RECT 16.900 72.800 17.800 73.100 ;
        RECT 19.000 73.000 21.000 73.100 ;
        RECT 16.900 71.100 17.300 72.800 ;
        RECT 19.000 71.100 19.400 73.000 ;
        RECT 20.600 71.100 21.000 73.000 ;
        RECT 21.400 71.100 21.800 73.100 ;
        RECT 22.200 73.000 24.200 73.100 ;
        RECT 22.200 71.100 22.600 73.000 ;
        RECT 23.800 71.100 24.200 73.000 ;
        RECT 24.600 71.100 25.000 73.100 ;
        RECT 25.700 72.800 26.600 73.100 ;
        RECT 25.700 71.100 26.100 72.800 ;
        RECT 27.800 72.400 28.200 73.200 ;
        RECT 28.600 71.100 29.000 75.800 ;
        RECT 29.400 74.800 29.800 75.200 ;
        RECT 29.400 74.200 29.700 74.800 ;
        RECT 30.400 74.200 30.700 75.900 ;
        RECT 33.400 75.800 34.400 76.200 ;
        RECT 34.700 75.900 35.400 76.200 ;
        RECT 35.000 75.800 35.400 75.900 ;
        RECT 31.000 75.100 31.400 75.200 ;
        RECT 33.400 75.100 33.800 75.200 ;
        RECT 31.000 74.800 33.800 75.100 ;
        RECT 31.000 74.400 31.400 74.800 ;
        RECT 33.400 74.400 33.800 74.800 ;
        RECT 34.100 74.200 34.400 75.800 ;
        RECT 29.400 73.800 30.700 74.200 ;
        RECT 31.800 74.100 32.200 74.200 ;
        RECT 32.600 74.100 33.000 74.200 ;
        RECT 31.400 73.800 33.400 74.100 ;
        RECT 34.100 73.800 35.400 74.200 ;
        RECT 29.500 73.100 29.800 73.800 ;
        RECT 31.400 73.600 31.800 73.800 ;
        RECT 33.000 73.600 33.400 73.800 ;
        RECT 30.300 73.100 32.100 73.300 ;
        RECT 32.700 73.100 34.500 73.300 ;
        RECT 35.000 73.100 35.300 73.800 ;
        RECT 36.600 73.100 37.000 79.900 ;
        RECT 38.200 75.900 38.600 79.900 ;
        RECT 39.000 76.200 39.400 79.900 ;
        RECT 40.600 76.200 41.000 79.900 ;
        RECT 41.400 77.900 41.800 79.900 ;
        RECT 41.500 77.800 41.800 77.900 ;
        RECT 43.000 77.800 43.400 79.900 ;
        RECT 41.500 77.500 43.300 77.800 ;
        RECT 41.500 76.200 41.800 77.500 ;
        RECT 42.200 76.400 42.600 77.200 ;
        RECT 39.000 75.900 41.000 76.200 ;
        RECT 38.300 75.200 38.600 75.900 ;
        RECT 41.400 75.800 41.800 76.200 ;
        RECT 44.600 75.900 45.000 79.900 ;
        RECT 45.400 76.200 45.800 79.900 ;
        RECT 47.000 76.200 47.400 79.900 ;
        RECT 50.200 77.900 50.600 79.900 ;
        RECT 50.300 77.800 50.600 77.900 ;
        RECT 51.800 77.900 52.200 79.900 ;
        RECT 51.800 77.800 52.100 77.900 ;
        RECT 50.300 77.500 52.100 77.800 ;
        RECT 51.000 76.400 51.400 77.200 ;
        RECT 51.800 76.200 52.100 77.500 ;
        RECT 45.400 75.900 47.400 76.200 ;
        RECT 38.200 74.900 39.400 75.200 ;
        RECT 38.200 74.800 38.600 74.900 ;
        RECT 38.200 74.100 38.600 74.200 ;
        RECT 39.100 74.100 39.400 74.900 ;
        RECT 38.200 73.800 39.400 74.100 ;
        RECT 41.500 74.200 41.800 75.800 ;
        RECT 44.700 75.200 45.000 75.900 ;
        RECT 49.400 75.400 49.800 76.200 ;
        RECT 51.800 75.800 52.200 76.200 ;
        RECT 44.600 74.900 45.800 75.200 ;
        RECT 44.600 74.800 45.000 74.900 ;
        RECT 41.500 74.100 42.300 74.200 ;
        RECT 41.500 73.900 42.400 74.100 ;
        RECT 29.400 71.100 29.800 73.100 ;
        RECT 30.200 73.000 32.200 73.100 ;
        RECT 30.200 71.100 30.600 73.000 ;
        RECT 31.800 71.100 32.200 73.000 ;
        RECT 32.600 73.000 34.600 73.100 ;
        RECT 32.600 71.100 33.000 73.000 ;
        RECT 34.200 71.100 34.600 73.000 ;
        RECT 35.000 71.100 35.400 73.100 ;
        RECT 36.100 72.800 37.000 73.100 ;
        RECT 38.200 72.800 38.600 73.200 ;
        RECT 39.100 73.100 39.400 73.800 ;
        RECT 36.100 72.200 36.500 72.800 ;
        RECT 38.300 72.400 38.700 72.800 ;
        RECT 35.800 71.800 36.500 72.200 ;
        RECT 36.100 71.100 36.500 71.800 ;
        RECT 39.000 71.100 39.400 73.100 ;
        RECT 42.000 71.100 42.400 73.900 ;
        RECT 45.500 73.200 45.800 74.900 ;
        RECT 50.200 74.800 51.000 75.200 ;
        RECT 51.800 74.200 52.100 75.800 ;
        RECT 51.300 74.100 52.100 74.200 ;
        RECT 44.600 72.800 45.000 73.200 ;
        RECT 44.700 72.400 45.100 72.800 ;
        RECT 45.400 71.100 45.800 73.200 ;
        RECT 51.200 73.900 52.100 74.100 ;
        RECT 51.200 71.100 51.600 73.900 ;
        RECT 52.600 71.100 53.000 79.900 ;
        RECT 55.000 77.900 55.400 79.900 ;
        RECT 55.100 77.800 55.400 77.900 ;
        RECT 56.600 77.900 57.000 79.900 ;
        RECT 56.600 77.800 56.900 77.900 ;
        RECT 58.200 77.800 58.600 79.900 ;
        RECT 59.800 77.900 60.200 79.900 ;
        RECT 60.900 79.200 61.300 79.900 ;
        RECT 60.600 78.800 61.300 79.200 ;
        RECT 59.800 77.800 60.100 77.900 ;
        RECT 55.100 77.500 56.900 77.800 ;
        RECT 58.300 77.500 60.100 77.800 ;
        RECT 55.800 76.400 56.200 77.200 ;
        RECT 56.600 76.200 56.900 77.500 ;
        RECT 59.000 76.400 59.400 77.200 ;
        RECT 59.800 76.200 60.100 77.500 ;
        RECT 60.900 76.300 61.300 78.800 ;
        RECT 64.100 79.200 64.500 79.900 ;
        RECT 67.500 79.200 67.900 79.900 ;
        RECT 70.700 79.200 71.100 79.900 ;
        RECT 73.100 79.200 73.500 79.900 ;
        RECT 64.100 78.800 65.000 79.200 ;
        RECT 67.000 78.800 67.900 79.200 ;
        RECT 70.200 78.800 71.100 79.200 ;
        RECT 72.600 78.800 73.500 79.200 ;
        RECT 63.400 76.800 63.800 77.200 ;
        RECT 53.400 76.100 53.800 76.200 ;
        RECT 54.200 76.100 54.600 76.200 ;
        RECT 53.400 75.800 54.600 76.100 ;
        RECT 54.200 75.400 54.600 75.800 ;
        RECT 56.600 75.800 57.000 76.200 ;
        RECT 59.800 75.800 60.200 76.200 ;
        RECT 60.900 75.900 61.800 76.300 ;
        RECT 63.400 76.200 63.700 76.800 ;
        RECT 64.100 76.200 64.500 78.800 ;
        RECT 63.000 75.900 63.700 76.200 ;
        RECT 64.000 75.900 64.500 76.200 ;
        RECT 67.500 76.200 67.900 78.800 ;
        RECT 68.200 76.800 68.600 77.200 ;
        RECT 68.300 76.200 68.600 76.800 ;
        RECT 70.700 76.300 71.100 78.800 ;
        RECT 67.500 75.900 68.000 76.200 ;
        RECT 68.300 75.900 69.000 76.200 ;
        RECT 70.200 75.900 71.100 76.300 ;
        RECT 73.100 76.200 73.500 78.800 ;
        RECT 73.800 76.800 74.200 77.200 ;
        RECT 73.900 76.200 74.200 76.800 ;
        RECT 75.800 77.100 76.200 79.900 ;
        RECT 76.600 77.100 77.000 77.200 ;
        RECT 75.800 76.800 77.000 77.100 ;
        RECT 73.100 75.900 73.600 76.200 ;
        RECT 73.900 75.900 74.600 76.200 ;
        RECT 55.000 74.800 55.800 75.200 ;
        RECT 56.600 74.200 56.900 75.800 ;
        RECT 59.800 74.200 60.100 75.800 ;
        RECT 60.600 74.800 61.000 75.600 ;
        RECT 56.100 74.100 56.900 74.200 ;
        RECT 59.300 74.100 60.100 74.200 ;
        RECT 56.000 73.900 56.900 74.100 ;
        RECT 59.200 73.900 60.100 74.100 ;
        RECT 61.400 74.200 61.700 75.900 ;
        RECT 63.000 75.800 63.400 75.900 ;
        RECT 64.000 74.200 64.300 75.900 ;
        RECT 64.600 75.100 65.000 75.200 ;
        RECT 67.000 75.100 67.400 75.200 ;
        RECT 64.600 74.800 67.400 75.100 ;
        RECT 64.600 74.400 65.000 74.800 ;
        RECT 67.000 74.400 67.400 74.800 ;
        RECT 67.700 74.200 68.000 75.900 ;
        RECT 68.600 75.800 69.000 75.900 ;
        RECT 70.300 74.200 70.600 75.900 ;
        RECT 71.000 74.800 71.400 75.600 ;
        RECT 72.600 74.400 73.000 75.200 ;
        RECT 73.300 74.200 73.600 75.900 ;
        RECT 74.200 75.800 74.600 75.900 ;
        RECT 53.400 72.400 53.800 73.200 ;
        RECT 56.000 71.100 56.400 73.900 ;
        RECT 59.200 71.100 59.600 73.900 ;
        RECT 61.400 73.800 61.800 74.200 ;
        RECT 63.000 73.800 64.300 74.200 ;
        RECT 65.400 74.100 65.800 74.200 ;
        RECT 66.200 74.100 66.600 74.200 ;
        RECT 65.000 73.800 67.000 74.100 ;
        RECT 67.700 73.800 69.000 74.200 ;
        RECT 70.200 73.800 70.600 74.200 ;
        RECT 71.800 74.100 72.200 74.200 ;
        RECT 71.800 73.800 72.600 74.100 ;
        RECT 73.300 73.800 74.600 74.200 ;
        RECT 61.400 72.100 61.700 73.800 ;
        RECT 62.200 72.400 62.600 73.200 ;
        RECT 63.100 73.100 63.400 73.800 ;
        RECT 65.000 73.600 65.400 73.800 ;
        RECT 66.600 73.600 67.000 73.800 ;
        RECT 63.900 73.100 65.700 73.300 ;
        RECT 66.300 73.100 68.100 73.300 ;
        RECT 68.600 73.100 68.900 73.800 ;
        RECT 61.400 71.100 61.800 72.100 ;
        RECT 63.000 71.100 63.400 73.100 ;
        RECT 63.800 73.000 65.800 73.100 ;
        RECT 63.800 71.100 64.200 73.000 ;
        RECT 65.400 71.100 65.800 73.000 ;
        RECT 66.200 73.000 68.200 73.100 ;
        RECT 66.200 71.100 66.600 73.000 ;
        RECT 67.800 71.100 68.200 73.000 ;
        RECT 68.600 71.100 69.000 73.100 ;
        RECT 69.400 72.400 69.800 73.200 ;
        RECT 70.300 72.100 70.600 73.800 ;
        RECT 72.200 73.600 72.600 73.800 ;
        RECT 71.900 73.100 73.700 73.300 ;
        RECT 74.200 73.100 74.500 73.800 ;
        RECT 75.000 73.400 75.400 74.200 ;
        RECT 70.200 71.100 70.600 72.100 ;
        RECT 71.800 73.000 73.800 73.100 ;
        RECT 71.800 71.100 72.200 73.000 ;
        RECT 73.400 71.100 73.800 73.000 ;
        RECT 74.200 71.100 74.600 73.100 ;
        RECT 75.800 71.100 76.200 76.800 ;
        RECT 76.600 73.400 77.000 74.200 ;
        RECT 77.400 73.100 77.800 79.900 ;
        RECT 77.400 72.800 78.300 73.100 ;
        RECT 77.900 72.200 78.300 72.800 ;
        RECT 77.900 71.800 78.600 72.200 ;
        RECT 77.900 71.100 78.300 71.800 ;
        RECT 79.800 71.100 80.200 79.900 ;
        RECT 82.200 75.100 82.600 79.900 ;
        RECT 85.100 76.200 85.500 79.900 ;
        RECT 87.300 79.200 87.700 79.900 ;
        RECT 87.300 78.800 88.200 79.200 ;
        RECT 85.800 76.800 86.200 77.200 ;
        RECT 85.900 76.200 86.200 76.800 ;
        RECT 87.300 76.300 87.700 78.800 ;
        RECT 85.100 75.900 85.600 76.200 ;
        RECT 85.900 75.900 86.600 76.200 ;
        RECT 87.300 75.900 88.200 76.300 ;
        RECT 90.700 76.200 91.100 79.900 ;
        RECT 91.400 76.800 91.800 77.200 ;
        RECT 91.500 76.200 91.800 76.800 ;
        RECT 90.700 75.900 91.200 76.200 ;
        RECT 91.500 75.900 92.200 76.200 ;
        RECT 84.600 75.100 85.000 75.200 ;
        RECT 80.600 74.800 82.600 75.100 ;
        RECT 80.600 74.200 80.900 74.800 ;
        RECT 80.600 73.800 81.000 74.200 ;
        RECT 81.400 73.400 81.800 74.200 ;
        RECT 82.200 73.100 82.600 74.800 ;
        RECT 83.000 74.800 85.000 75.100 ;
        RECT 83.000 74.200 83.300 74.800 ;
        RECT 84.600 74.400 85.000 74.800 ;
        RECT 85.300 74.200 85.600 75.900 ;
        RECT 86.200 75.800 86.600 75.900 ;
        RECT 86.200 75.100 86.600 75.200 ;
        RECT 87.000 75.100 87.400 75.600 ;
        RECT 86.200 74.800 87.400 75.100 ;
        RECT 87.800 74.200 88.100 75.900 ;
        RECT 90.200 74.400 90.600 75.200 ;
        RECT 90.900 74.200 91.200 75.900 ;
        RECT 91.800 75.800 92.200 75.900 ;
        RECT 83.000 73.800 83.400 74.200 ;
        RECT 83.800 74.100 84.200 74.200 ;
        RECT 85.300 74.100 86.600 74.200 ;
        RECT 87.000 74.100 87.400 74.200 ;
        RECT 83.800 73.800 84.600 74.100 ;
        RECT 85.300 73.800 87.400 74.100 ;
        RECT 87.800 73.800 88.200 74.200 ;
        RECT 89.400 74.100 89.800 74.200 ;
        RECT 89.400 73.800 90.200 74.100 ;
        RECT 90.900 73.800 92.200 74.200 ;
        RECT 84.200 73.600 84.600 73.800 ;
        RECT 83.900 73.100 85.700 73.300 ;
        RECT 86.200 73.100 86.500 73.800 ;
        RECT 82.200 72.800 83.100 73.100 ;
        RECT 82.700 71.100 83.100 72.800 ;
        RECT 83.800 73.000 85.800 73.100 ;
        RECT 83.800 71.100 84.200 73.000 ;
        RECT 85.400 71.100 85.800 73.000 ;
        RECT 86.200 71.100 86.600 73.100 ;
        RECT 87.800 72.100 88.100 73.800 ;
        RECT 89.800 73.600 90.200 73.800 ;
        RECT 88.600 72.400 89.000 73.200 ;
        RECT 89.500 73.100 91.300 73.300 ;
        RECT 91.800 73.100 92.100 73.800 ;
        RECT 92.600 73.400 93.000 74.200 ;
        RECT 93.400 73.200 93.800 79.900 ;
        RECT 95.800 77.900 96.200 79.900 ;
        RECT 94.200 75.800 94.600 76.600 ;
        RECT 95.900 75.800 96.200 77.900 ;
        RECT 97.400 75.900 97.800 79.900 ;
        RECT 98.200 79.600 100.200 79.900 ;
        RECT 98.200 75.900 98.600 79.600 ;
        RECT 99.000 75.900 99.400 79.300 ;
        RECT 99.800 76.200 100.200 79.600 ;
        RECT 101.400 76.200 101.800 79.900 ;
        RECT 99.800 75.900 101.800 76.200 ;
        RECT 95.900 75.500 97.100 75.800 ;
        RECT 95.800 74.800 96.200 75.200 ;
        RECT 94.200 73.800 94.600 74.200 ;
        RECT 95.000 73.800 95.400 74.600 ;
        RECT 95.900 74.400 96.200 74.800 ;
        RECT 95.900 74.100 96.400 74.400 ;
        RECT 96.000 74.000 96.400 74.100 ;
        RECT 96.800 73.800 97.100 75.500 ;
        RECT 97.500 75.200 97.800 75.900 ;
        RECT 99.100 75.600 99.400 75.900 ;
        RECT 97.400 75.100 97.800 75.200 ;
        RECT 98.200 75.100 98.600 75.600 ;
        RECT 99.100 75.300 100.100 75.600 ;
        RECT 97.400 74.800 98.600 75.100 ;
        RECT 99.800 75.200 100.100 75.300 ;
        RECT 101.000 75.200 101.400 75.400 ;
        RECT 99.800 74.800 100.200 75.200 ;
        RECT 101.000 74.900 101.800 75.200 ;
        RECT 101.400 74.800 101.800 74.900 ;
        RECT 94.200 73.200 94.500 73.800 ;
        RECT 96.800 73.700 97.200 73.800 ;
        RECT 95.700 73.500 97.200 73.700 ;
        RECT 89.400 73.000 91.400 73.100 ;
        RECT 87.800 71.100 88.200 72.100 ;
        RECT 89.400 71.100 89.800 73.000 ;
        RECT 91.000 71.100 91.400 73.000 ;
        RECT 91.800 71.100 92.200 73.100 ;
        RECT 93.400 72.800 94.500 73.200 ;
        RECT 95.100 73.400 97.200 73.500 ;
        RECT 95.100 73.200 96.000 73.400 ;
        RECT 95.100 73.100 95.400 73.200 ;
        RECT 97.500 73.100 97.800 74.800 ;
        RECT 99.100 74.400 99.500 74.800 ;
        RECT 99.100 74.200 99.400 74.400 ;
        RECT 99.000 73.800 99.400 74.200 ;
        RECT 99.800 73.100 100.100 74.800 ;
        RECT 100.600 74.100 101.000 74.600 ;
        RECT 103.000 74.100 103.400 74.200 ;
        RECT 100.600 73.800 103.400 74.100 ;
        RECT 93.900 71.100 94.300 72.800 ;
        RECT 95.000 71.100 95.400 73.100 ;
        RECT 97.100 72.600 97.800 73.100 ;
        RECT 97.100 71.100 97.500 72.600 ;
        RECT 99.500 72.200 100.300 73.100 ;
        RECT 99.000 71.800 100.300 72.200 ;
        RECT 99.500 71.100 100.300 71.800 ;
        RECT 103.800 71.100 104.200 79.900 ;
        RECT 105.400 75.900 105.800 79.900 ;
        RECT 106.200 76.200 106.600 79.900 ;
        RECT 107.800 76.200 108.200 79.900 ;
        RECT 106.200 75.900 108.200 76.200 ;
        RECT 108.600 76.200 109.000 79.900 ;
        RECT 110.200 76.200 110.600 79.900 ;
        RECT 108.600 75.900 110.600 76.200 ;
        RECT 111.000 75.900 111.400 79.900 ;
        RECT 111.800 75.900 112.200 79.900 ;
        RECT 113.400 77.900 113.800 79.900 ;
        RECT 105.500 75.200 105.800 75.900 ;
        RECT 107.400 75.200 107.800 75.400 ;
        RECT 111.000 75.200 111.300 75.900 ;
        RECT 111.800 75.200 112.100 75.900 ;
        RECT 113.400 75.800 113.700 77.900 ;
        RECT 115.300 76.300 115.700 79.900 ;
        RECT 118.500 79.200 118.900 79.900 ;
        RECT 118.500 78.800 119.400 79.200 ;
        RECT 117.800 76.800 118.200 77.200 ;
        RECT 115.300 75.900 116.200 76.300 ;
        RECT 117.800 76.200 118.100 76.800 ;
        RECT 118.500 76.200 118.900 78.800 ;
        RECT 117.400 75.900 118.100 76.200 ;
        RECT 118.400 75.900 118.900 76.200 ;
        RECT 112.500 75.500 113.700 75.800 ;
        RECT 105.400 74.900 106.600 75.200 ;
        RECT 107.400 74.900 108.200 75.200 ;
        RECT 105.400 74.800 105.800 74.900 ;
        RECT 104.600 72.400 105.000 73.200 ;
        RECT 105.400 72.800 105.800 73.200 ;
        RECT 106.300 73.100 106.600 74.900 ;
        RECT 107.800 74.800 108.200 74.900 ;
        RECT 110.200 74.900 111.400 75.200 ;
        RECT 107.000 73.800 107.400 74.600 ;
        RECT 108.600 74.100 109.000 74.200 ;
        RECT 109.400 74.100 109.800 74.600 ;
        RECT 108.600 73.800 109.800 74.100 ;
        RECT 105.500 72.400 105.900 72.800 ;
        RECT 106.200 71.100 106.600 73.100 ;
        RECT 110.200 73.100 110.500 74.900 ;
        RECT 111.000 74.800 111.400 74.900 ;
        RECT 111.800 74.800 112.200 75.200 ;
        RECT 110.200 71.100 110.600 73.100 ;
        RECT 111.000 72.800 111.400 73.200 ;
        RECT 111.800 73.100 112.100 74.800 ;
        RECT 112.500 73.800 112.800 75.500 ;
        RECT 113.400 74.800 113.800 75.200 ;
        RECT 115.000 74.800 115.400 75.600 ;
        RECT 115.800 75.100 116.100 75.900 ;
        RECT 117.400 75.800 117.800 75.900 ;
        RECT 117.400 75.100 117.700 75.800 ;
        RECT 115.800 74.800 117.700 75.100 ;
        RECT 113.400 74.400 113.700 74.800 ;
        RECT 113.200 74.100 113.700 74.400 ;
        RECT 113.200 74.000 113.600 74.100 ;
        RECT 114.200 73.800 114.600 74.600 ;
        RECT 115.800 74.200 116.100 74.800 ;
        RECT 118.400 74.200 118.700 75.900 ;
        RECT 120.600 75.800 121.000 76.600 ;
        RECT 119.000 74.400 119.400 75.200 ;
        RECT 119.800 75.100 120.200 75.200 ;
        RECT 120.600 75.100 120.900 75.800 ;
        RECT 119.800 74.800 120.900 75.100 ;
        RECT 115.800 73.800 116.200 74.200 ;
        RECT 117.400 73.800 118.700 74.200 ;
        RECT 119.800 74.100 120.200 74.200 ;
        RECT 121.400 74.100 121.800 79.900 ;
        RECT 123.000 75.900 123.400 79.900 ;
        RECT 123.800 76.200 124.200 79.900 ;
        RECT 125.400 76.200 125.800 79.900 ;
        RECT 127.000 77.900 127.400 79.900 ;
        RECT 123.800 75.900 125.800 76.200 ;
        RECT 123.100 75.200 123.400 75.900 ;
        RECT 127.100 75.800 127.400 77.900 ;
        RECT 128.600 75.900 129.000 79.900 ;
        RECT 129.700 76.300 130.100 79.900 ;
        RECT 129.700 75.900 130.600 76.300 ;
        RECT 127.100 75.500 128.300 75.800 ;
        RECT 125.000 75.200 125.400 75.400 ;
        RECT 123.000 74.900 124.200 75.200 ;
        RECT 125.000 74.900 125.800 75.200 ;
        RECT 123.000 74.800 123.400 74.900 ;
        RECT 119.400 73.800 121.800 74.100 ;
        RECT 112.400 73.700 112.800 73.800 ;
        RECT 112.400 73.500 113.900 73.700 ;
        RECT 112.400 73.400 114.500 73.500 ;
        RECT 113.600 73.200 114.500 73.400 ;
        RECT 114.200 73.100 114.500 73.200 ;
        RECT 110.900 72.400 111.300 72.800 ;
        RECT 111.800 72.600 112.500 73.100 ;
        RECT 112.100 72.200 112.500 72.600 ;
        RECT 111.800 71.800 112.500 72.200 ;
        RECT 112.100 71.100 112.500 71.800 ;
        RECT 114.200 71.100 114.600 73.100 ;
        RECT 115.800 72.100 116.100 73.800 ;
        RECT 116.600 72.400 117.000 73.200 ;
        RECT 117.500 73.100 117.800 73.800 ;
        RECT 119.400 73.600 119.800 73.800 ;
        RECT 118.300 73.100 120.100 73.300 ;
        RECT 121.400 73.100 121.800 73.800 ;
        RECT 122.200 73.400 122.600 74.200 ;
        RECT 115.800 71.100 116.200 72.100 ;
        RECT 117.400 71.100 117.800 73.100 ;
        RECT 118.200 73.000 120.200 73.100 ;
        RECT 118.200 71.100 118.600 73.000 ;
        RECT 119.800 71.100 120.200 73.000 ;
        RECT 120.900 72.800 121.800 73.100 ;
        RECT 123.000 72.800 123.400 73.200 ;
        RECT 123.900 73.100 124.200 74.900 ;
        RECT 125.400 74.800 125.800 74.900 ;
        RECT 127.000 74.800 127.400 75.200 ;
        RECT 124.600 73.800 125.000 74.600 ;
        RECT 126.200 73.800 126.600 74.600 ;
        RECT 127.100 74.400 127.400 74.800 ;
        RECT 127.100 74.100 127.600 74.400 ;
        RECT 127.200 74.000 127.600 74.100 ;
        RECT 128.000 73.800 128.300 75.500 ;
        RECT 128.700 75.200 129.000 75.900 ;
        RECT 128.600 74.800 129.000 75.200 ;
        RECT 129.400 74.800 129.800 75.600 ;
        RECT 128.000 73.700 128.400 73.800 ;
        RECT 126.900 73.500 128.400 73.700 ;
        RECT 126.300 73.400 128.400 73.500 ;
        RECT 126.300 73.200 127.200 73.400 ;
        RECT 126.300 73.100 126.600 73.200 ;
        RECT 128.700 73.100 129.000 74.800 ;
        RECT 130.200 74.200 130.500 75.900 ;
        RECT 129.400 74.100 129.800 74.200 ;
        RECT 130.200 74.100 130.600 74.200 ;
        RECT 131.800 74.100 132.200 74.200 ;
        RECT 129.400 73.800 130.600 74.100 ;
        RECT 131.000 73.800 132.200 74.100 ;
        RECT 120.900 71.100 121.300 72.800 ;
        RECT 123.100 72.400 123.500 72.800 ;
        RECT 123.800 71.100 124.200 73.100 ;
        RECT 126.200 71.100 126.600 73.100 ;
        RECT 128.300 72.600 129.000 73.100 ;
        RECT 128.300 71.100 128.700 72.600 ;
        RECT 130.200 72.100 130.500 73.800 ;
        RECT 131.000 73.200 131.300 73.800 ;
        RECT 131.800 73.400 132.200 73.800 ;
        RECT 131.000 72.400 131.400 73.200 ;
        RECT 130.200 71.100 130.600 72.100 ;
        RECT 132.600 71.100 133.000 79.900 ;
        RECT 134.700 76.200 135.100 79.900 ;
        RECT 137.900 77.200 138.300 79.900 ;
        RECT 140.900 79.200 141.300 79.900 ;
        RECT 140.900 78.800 141.800 79.200 ;
        RECT 135.400 76.800 135.800 77.200 ;
        RECT 137.400 76.800 138.300 77.200 ;
        RECT 138.600 76.800 139.000 77.200 ;
        RECT 135.500 76.200 135.800 76.800 ;
        RECT 137.900 76.200 138.300 76.800 ;
        RECT 138.700 76.200 139.000 76.800 ;
        RECT 140.900 76.200 141.300 78.800 ;
        RECT 134.700 75.900 135.200 76.200 ;
        RECT 135.500 75.900 136.200 76.200 ;
        RECT 137.900 75.900 138.400 76.200 ;
        RECT 138.700 75.900 139.400 76.200 ;
        RECT 134.200 74.400 134.600 75.200 ;
        RECT 134.900 74.200 135.200 75.900 ;
        RECT 135.800 75.800 136.200 75.900 ;
        RECT 135.800 74.800 136.200 75.200 ;
        RECT 135.800 74.200 136.100 74.800 ;
        RECT 137.400 74.400 137.800 75.200 ;
        RECT 138.100 74.200 138.400 75.900 ;
        RECT 139.000 75.800 139.400 75.900 ;
        RECT 140.800 75.900 141.300 76.200 ;
        RECT 140.800 74.200 141.100 75.900 ;
        RECT 143.000 75.600 143.400 79.900 ;
        RECT 145.100 76.200 145.500 79.900 ;
        RECT 145.100 75.900 145.800 76.200 ;
        RECT 143.000 75.400 145.000 75.600 ;
        RECT 143.000 75.300 145.100 75.400 ;
        RECT 141.400 74.400 141.800 75.200 ;
        RECT 144.700 75.000 145.100 75.300 ;
        RECT 145.500 75.200 145.800 75.900 ;
        RECT 144.000 74.200 144.400 74.600 ;
        RECT 133.400 74.100 133.800 74.200 ;
        RECT 133.400 73.800 134.200 74.100 ;
        RECT 134.900 73.800 136.200 74.200 ;
        RECT 136.600 74.100 137.000 74.200 ;
        RECT 136.600 73.800 137.400 74.100 ;
        RECT 138.100 73.800 139.400 74.200 ;
        RECT 139.800 73.800 141.100 74.200 ;
        RECT 142.200 74.100 142.600 74.200 ;
        RECT 141.800 73.800 142.600 74.100 ;
        RECT 143.800 73.800 144.300 74.200 ;
        RECT 133.800 73.600 134.200 73.800 ;
        RECT 133.500 73.100 135.300 73.300 ;
        RECT 135.800 73.100 136.100 73.800 ;
        RECT 137.000 73.600 137.400 73.800 ;
        RECT 136.700 73.100 138.500 73.300 ;
        RECT 139.000 73.100 139.300 73.800 ;
        RECT 139.900 73.100 140.200 73.800 ;
        RECT 141.800 73.600 142.200 73.800 ;
        RECT 144.800 73.500 145.100 75.000 ;
        RECT 145.400 74.800 145.800 75.200 ;
        RECT 140.700 73.100 142.500 73.300 ;
        RECT 143.900 73.200 145.100 73.500 ;
        RECT 133.400 73.000 135.400 73.100 ;
        RECT 133.400 71.100 133.800 73.000 ;
        RECT 135.000 71.100 135.400 73.000 ;
        RECT 135.800 71.100 136.200 73.100 ;
        RECT 136.600 73.000 138.600 73.100 ;
        RECT 136.600 71.100 137.000 73.000 ;
        RECT 138.200 71.100 138.600 73.000 ;
        RECT 139.000 71.100 139.400 73.100 ;
        RECT 139.800 71.100 140.200 73.100 ;
        RECT 140.600 73.000 142.600 73.100 ;
        RECT 140.600 71.100 141.000 73.000 ;
        RECT 142.200 71.100 142.600 73.000 ;
        RECT 143.000 72.400 143.400 73.200 ;
        RECT 143.900 72.100 144.200 73.200 ;
        RECT 145.500 73.100 145.800 74.800 ;
        RECT 143.800 71.100 144.200 72.100 ;
        RECT 145.400 71.100 145.800 73.100 ;
        RECT 146.200 71.100 146.600 79.900 ;
        RECT 147.000 74.100 147.400 74.200 ;
        RECT 147.800 74.100 148.200 74.200 ;
        RECT 147.000 73.800 148.200 74.100 ;
        RECT 147.000 73.400 147.400 73.800 ;
        RECT 147.800 73.400 148.200 73.800 ;
        RECT 148.600 73.100 149.000 79.900 ;
        RECT 149.400 76.100 149.800 76.600 ;
        RECT 150.200 76.100 150.600 76.200 ;
        RECT 149.400 75.800 150.600 76.100 ;
        RECT 148.600 72.800 149.500 73.100 ;
        RECT 149.100 72.200 149.500 72.800 ;
        RECT 148.600 71.800 149.500 72.200 ;
        RECT 149.100 71.100 149.500 71.800 ;
        RECT 2.200 67.900 2.600 69.900 ;
        RECT 4.600 68.800 5.000 69.900 ;
        RECT 2.900 68.200 3.300 68.600 ;
        RECT 1.400 66.400 1.800 67.200 ;
        RECT 2.200 67.100 2.500 67.900 ;
        RECT 3.000 67.800 3.400 68.200 ;
        RECT 3.800 67.800 4.200 68.600 ;
        RECT 3.800 67.100 4.100 67.800 ;
        RECT 4.700 67.200 5.000 68.800 ;
        RECT 6.300 68.200 6.700 68.600 ;
        RECT 5.400 68.100 5.800 68.200 ;
        RECT 6.200 68.100 6.600 68.200 ;
        RECT 5.400 67.800 6.600 68.100 ;
        RECT 7.000 67.900 7.400 69.900 ;
        RECT 11.200 69.200 11.600 69.900 ;
        RECT 13.200 69.200 13.600 69.900 ;
        RECT 11.000 68.800 11.600 69.200 ;
        RECT 12.600 68.800 13.600 69.200 ;
        RECT 16.600 69.100 17.000 69.200 ;
        RECT 17.600 69.100 18.000 69.900 ;
        RECT 16.600 68.800 18.000 69.100 ;
        RECT 2.200 66.800 4.100 67.100 ;
        RECT 4.600 66.800 5.000 67.200 ;
        RECT 0.600 66.100 1.000 66.200 ;
        RECT 2.200 66.100 2.500 66.800 ;
        RECT 3.000 66.100 3.400 66.200 ;
        RECT 0.600 65.800 1.400 66.100 ;
        RECT 2.200 65.800 3.400 66.100 ;
        RECT 1.000 65.600 1.400 65.800 ;
        RECT 3.000 65.100 3.300 65.800 ;
        RECT 4.700 65.100 5.000 66.800 ;
        RECT 5.400 66.100 5.800 66.200 ;
        RECT 6.200 66.100 6.600 66.200 ;
        RECT 7.100 66.100 7.400 67.900 ;
        RECT 7.800 66.400 8.200 67.200 ;
        RECT 11.200 67.100 11.600 68.800 ;
        RECT 13.200 67.100 13.600 68.800 ;
        RECT 11.200 66.900 12.100 67.100 ;
        RECT 11.300 66.800 12.100 66.900 ;
        RECT 8.600 66.100 9.000 66.200 ;
        RECT 5.400 65.800 7.400 66.100 ;
        RECT 8.200 65.800 9.000 66.100 ;
        RECT 10.200 65.800 11.000 66.200 ;
        RECT 5.400 65.400 5.800 65.800 ;
        RECT 6.300 65.100 6.600 65.800 ;
        RECT 8.200 65.600 8.600 65.800 ;
        RECT 0.600 64.800 2.600 65.100 ;
        RECT 0.600 61.100 1.000 64.800 ;
        RECT 2.200 61.100 2.600 64.800 ;
        RECT 3.000 61.100 3.400 65.100 ;
        RECT 4.600 64.700 5.500 65.100 ;
        RECT 5.100 61.100 5.500 64.700 ;
        RECT 6.200 61.100 6.600 65.100 ;
        RECT 7.000 64.800 9.000 65.100 ;
        RECT 9.400 64.800 9.800 65.600 ;
        RECT 11.800 65.200 12.100 66.800 ;
        RECT 12.700 66.900 13.600 67.100 ;
        RECT 17.600 67.100 18.000 68.800 ;
        RECT 19.300 68.400 19.700 69.900 ;
        RECT 19.000 67.900 19.700 68.400 ;
        RECT 21.400 67.900 21.800 69.900 ;
        RECT 23.000 68.800 23.400 69.900 ;
        RECT 24.600 69.600 26.600 69.900 ;
        RECT 17.600 66.900 18.500 67.100 ;
        RECT 12.700 66.800 13.500 66.900 ;
        RECT 17.700 66.800 18.500 66.900 ;
        RECT 12.700 65.200 13.000 66.800 ;
        RECT 13.800 65.800 14.600 66.200 ;
        RECT 16.600 65.800 17.400 66.200 ;
        RECT 11.800 64.800 12.200 65.200 ;
        RECT 12.600 64.800 13.000 65.200 ;
        RECT 15.000 64.800 15.400 65.600 ;
        RECT 15.800 64.800 16.200 65.600 ;
        RECT 18.200 65.200 18.500 66.800 ;
        RECT 19.000 66.200 19.300 67.900 ;
        RECT 21.400 67.800 21.700 67.900 ;
        RECT 20.800 67.600 21.700 67.800 ;
        RECT 19.600 67.500 21.700 67.600 ;
        RECT 19.600 67.300 21.100 67.500 ;
        RECT 19.600 67.200 20.000 67.300 ;
        RECT 23.000 67.200 23.300 68.800 ;
        RECT 23.800 67.800 24.200 68.600 ;
        RECT 24.600 67.900 25.000 69.600 ;
        RECT 25.400 67.900 25.800 69.300 ;
        RECT 26.200 68.000 26.600 69.600 ;
        RECT 27.800 68.000 28.200 69.900 ;
        RECT 28.900 68.200 29.300 69.900 ;
        RECT 31.100 68.200 31.500 68.600 ;
        RECT 26.200 67.900 28.200 68.000 ;
        RECT 25.400 67.200 25.700 67.900 ;
        RECT 26.300 67.700 28.100 67.900 ;
        RECT 28.600 67.800 29.800 68.200 ;
        RECT 31.000 67.800 31.400 68.200 ;
        RECT 31.800 67.900 32.200 69.900 ;
        RECT 34.500 69.200 34.900 69.900 ;
        RECT 36.900 69.200 37.300 69.900 ;
        RECT 34.200 68.800 34.900 69.200 ;
        RECT 36.600 68.800 37.300 69.200 ;
        RECT 34.500 68.200 34.900 68.800 ;
        RECT 36.900 68.200 37.300 68.800 ;
        RECT 34.500 67.900 35.400 68.200 ;
        RECT 36.900 67.900 37.800 68.200 ;
        RECT 39.000 67.900 39.400 69.900 ;
        RECT 39.800 68.000 40.200 69.900 ;
        RECT 41.400 68.000 41.800 69.900 ;
        RECT 39.800 67.900 41.800 68.000 ;
        RECT 42.200 68.000 42.600 69.900 ;
        RECT 43.800 68.000 44.200 69.900 ;
        RECT 42.200 67.900 44.200 68.000 ;
        RECT 44.600 67.900 45.000 69.900 ;
        RECT 45.400 67.900 45.800 69.900 ;
        RECT 46.200 68.000 46.600 69.900 ;
        RECT 47.800 68.000 48.200 69.900 ;
        RECT 46.200 67.900 48.200 68.000 ;
        RECT 50.200 68.000 50.600 69.900 ;
        RECT 51.800 68.000 52.200 69.900 ;
        RECT 50.200 67.900 52.200 68.000 ;
        RECT 52.600 67.900 53.000 69.900 ;
        RECT 53.700 69.200 54.100 69.900 ;
        RECT 53.400 68.800 54.100 69.200 ;
        RECT 53.700 68.200 54.100 68.800 ;
        RECT 53.700 67.900 54.600 68.200 ;
        RECT 55.800 68.000 56.200 69.900 ;
        RECT 57.400 69.600 59.400 69.900 ;
        RECT 57.400 68.000 57.800 69.600 ;
        RECT 55.800 67.900 57.800 68.000 ;
        RECT 58.200 67.900 58.600 69.300 ;
        RECT 59.000 67.900 59.400 69.600 ;
        RECT 61.100 68.200 61.900 69.900 ;
        RECT 63.900 68.200 64.300 68.600 ;
        RECT 60.600 67.900 61.900 68.200 ;
        RECT 27.400 67.200 27.800 67.400 ;
        RECT 28.600 67.200 28.900 67.800 ;
        RECT 19.000 65.800 19.400 66.200 ;
        RECT 18.200 64.800 18.600 65.200 ;
        RECT 19.000 65.100 19.300 65.800 ;
        RECT 19.700 65.500 20.000 67.200 ;
        RECT 20.400 66.900 20.800 67.000 ;
        RECT 20.400 66.600 20.900 66.900 ;
        RECT 20.600 66.200 20.900 66.600 ;
        RECT 21.400 66.400 21.800 67.200 ;
        RECT 23.000 66.800 23.400 67.200 ;
        RECT 23.800 66.800 24.200 67.200 ;
        RECT 20.600 65.800 21.000 66.200 ;
        RECT 19.700 65.200 20.900 65.500 ;
        RECT 22.200 65.400 22.600 66.200 ;
        RECT 7.000 61.100 7.400 64.800 ;
        RECT 8.600 61.100 9.000 64.800 ;
        RECT 11.000 63.800 11.400 64.600 ;
        RECT 11.800 63.500 12.100 64.800 ;
        RECT 10.300 63.200 12.100 63.500 ;
        RECT 10.300 63.100 10.600 63.200 ;
        RECT 10.200 61.100 10.600 63.100 ;
        RECT 11.800 63.100 12.100 63.200 ;
        RECT 12.700 63.500 13.000 64.800 ;
        RECT 13.400 64.100 13.800 64.600 ;
        RECT 16.600 64.100 17.000 64.200 ;
        RECT 17.400 64.100 17.800 64.600 ;
        RECT 13.400 63.800 17.800 64.100 ;
        RECT 18.200 63.500 18.500 64.800 ;
        RECT 12.700 63.200 14.500 63.500 ;
        RECT 12.700 63.100 13.000 63.200 ;
        RECT 11.800 61.100 12.200 63.100 ;
        RECT 12.600 61.100 13.000 63.100 ;
        RECT 14.200 63.100 14.500 63.200 ;
        RECT 16.700 63.200 18.500 63.500 ;
        RECT 16.700 63.100 17.000 63.200 ;
        RECT 14.200 61.100 14.600 63.100 ;
        RECT 16.600 61.100 17.000 63.100 ;
        RECT 18.200 63.100 18.500 63.200 ;
        RECT 18.200 61.100 18.600 63.100 ;
        RECT 19.000 61.100 19.400 65.100 ;
        RECT 20.600 63.100 20.900 65.200 ;
        RECT 23.000 65.100 23.300 66.800 ;
        RECT 23.800 66.100 24.100 66.800 ;
        RECT 24.600 66.100 25.000 67.200 ;
        RECT 25.400 66.900 26.600 67.200 ;
        RECT 27.400 66.900 28.200 67.200 ;
        RECT 26.200 66.800 26.600 66.900 ;
        RECT 27.800 66.800 28.200 66.900 ;
        RECT 28.600 66.800 29.000 67.200 ;
        RECT 23.800 65.800 25.000 66.100 ;
        RECT 25.400 65.800 25.800 66.600 ;
        RECT 26.300 65.100 26.600 66.800 ;
        RECT 27.000 65.800 27.400 66.600 ;
        RECT 22.500 64.700 23.400 65.100 ;
        RECT 20.600 61.100 21.000 63.100 ;
        RECT 22.500 61.100 22.900 64.700 ;
        RECT 25.900 63.200 26.900 65.100 ;
        RECT 25.400 62.800 26.900 63.200 ;
        RECT 25.900 61.100 26.900 62.800 ;
        RECT 29.400 61.100 29.800 67.800 ;
        RECT 31.000 66.100 31.400 66.200 ;
        RECT 31.900 66.100 32.200 67.900 ;
        RECT 31.000 65.800 32.200 66.100 ;
        RECT 31.100 65.100 31.400 65.800 ;
        RECT 31.000 61.100 31.400 65.100 ;
        RECT 31.800 64.800 33.800 65.100 ;
        RECT 31.800 61.100 32.200 64.800 ;
        RECT 33.400 61.100 33.800 64.800 ;
        RECT 35.000 61.100 35.400 67.900 ;
        RECT 37.400 61.100 37.800 67.900 ;
        RECT 39.100 67.200 39.400 67.900 ;
        RECT 39.900 67.700 41.700 67.900 ;
        RECT 42.300 67.700 44.100 67.900 ;
        RECT 41.000 67.200 41.400 67.400 ;
        RECT 42.600 67.200 43.000 67.400 ;
        RECT 44.600 67.200 44.900 67.900 ;
        RECT 45.500 67.200 45.800 67.900 ;
        RECT 46.300 67.700 48.100 67.900 ;
        RECT 50.300 67.700 52.100 67.900 ;
        RECT 47.400 67.200 47.800 67.400 ;
        RECT 50.600 67.200 51.000 67.400 ;
        RECT 52.600 67.200 52.900 67.900 ;
        RECT 39.000 66.800 40.300 67.200 ;
        RECT 41.000 67.100 41.800 67.200 ;
        RECT 42.200 67.100 43.000 67.200 ;
        RECT 41.000 66.900 43.000 67.100 ;
        RECT 41.400 66.800 42.600 66.900 ;
        RECT 43.700 66.800 45.000 67.200 ;
        RECT 45.400 66.800 46.700 67.200 ;
        RECT 47.400 67.100 48.200 67.200 ;
        RECT 50.200 67.100 51.000 67.200 ;
        RECT 47.400 66.900 51.000 67.100 ;
        RECT 47.800 66.800 50.600 66.900 ;
        RECT 51.700 66.800 53.000 67.200 ;
        RECT 39.000 65.100 39.400 65.200 ;
        RECT 40.000 65.100 40.300 66.800 ;
        RECT 40.600 66.100 41.000 66.600 ;
        RECT 43.000 66.100 43.400 66.600 ;
        RECT 40.600 65.800 43.400 66.100 ;
        RECT 43.700 65.100 44.000 66.800 ;
        RECT 44.600 65.100 45.000 65.200 ;
        RECT 45.400 65.100 45.800 65.200 ;
        RECT 46.400 65.100 46.700 66.800 ;
        RECT 47.000 66.100 47.400 66.600 ;
        RECT 51.000 66.100 51.400 66.600 ;
        RECT 47.000 65.800 51.400 66.100 ;
        RECT 51.700 65.100 52.000 66.800 ;
        RECT 52.600 65.100 53.000 65.200 ;
        RECT 39.000 64.800 39.700 65.100 ;
        RECT 40.000 64.800 40.500 65.100 ;
        RECT 39.400 64.200 39.700 64.800 ;
        RECT 39.400 63.800 39.800 64.200 ;
        RECT 40.100 61.100 40.500 64.800 ;
        RECT 43.500 64.800 44.000 65.100 ;
        RECT 44.300 64.800 46.100 65.100 ;
        RECT 46.400 64.800 46.900 65.100 ;
        RECT 43.500 61.100 43.900 64.800 ;
        RECT 44.300 64.200 44.600 64.800 ;
        RECT 44.200 63.800 44.600 64.200 ;
        RECT 45.800 64.200 46.100 64.800 ;
        RECT 45.800 63.800 46.200 64.200 ;
        RECT 46.500 61.100 46.900 64.800 ;
        RECT 51.500 64.800 52.000 65.100 ;
        RECT 52.300 64.800 53.000 65.100 ;
        RECT 51.500 61.100 51.900 64.800 ;
        RECT 52.300 64.200 52.600 64.800 ;
        RECT 52.200 63.800 52.600 64.200 ;
        RECT 54.200 61.100 54.600 67.900 ;
        RECT 55.900 67.700 57.700 67.900 ;
        RECT 56.200 67.200 56.600 67.400 ;
        RECT 58.300 67.200 58.600 67.900 ;
        RECT 60.600 67.800 61.700 67.900 ;
        RECT 63.800 67.800 64.200 68.200 ;
        RECT 64.600 67.900 65.000 69.900 ;
        RECT 55.800 66.900 56.600 67.200 ;
        RECT 57.400 66.900 58.600 67.200 ;
        RECT 59.000 67.100 59.400 67.200 ;
        RECT 59.800 67.100 60.200 67.200 ;
        RECT 55.800 66.800 56.200 66.900 ;
        RECT 57.400 66.800 57.800 66.900 ;
        RECT 59.000 66.800 60.200 67.100 ;
        RECT 60.600 66.800 61.000 67.200 ;
        RECT 56.600 65.800 57.000 66.600 ;
        RECT 57.400 65.100 57.700 66.800 ;
        RECT 58.200 65.800 58.600 66.600 ;
        RECT 59.000 66.400 59.400 66.800 ;
        RECT 60.700 66.600 61.000 66.800 ;
        RECT 60.700 66.200 61.100 66.600 ;
        RECT 61.400 66.200 61.700 67.800 ;
        RECT 61.400 65.800 61.800 66.200 ;
        RECT 63.000 66.100 63.400 66.200 ;
        RECT 62.600 65.800 63.400 66.100 ;
        RECT 63.800 66.100 64.200 66.200 ;
        RECT 64.700 66.100 65.000 67.900 ;
        RECT 68.600 67.900 69.000 69.900 ;
        RECT 71.500 69.200 71.900 69.900 ;
        RECT 71.000 68.800 71.900 69.200 ;
        RECT 69.300 68.200 69.700 68.600 ;
        RECT 71.500 68.200 71.900 68.800 ;
        RECT 65.400 66.400 65.800 67.200 ;
        RECT 63.800 65.800 65.000 66.100 ;
        RECT 67.000 66.100 67.400 66.200 ;
        RECT 68.600 66.100 68.900 67.900 ;
        RECT 69.400 67.800 69.800 68.200 ;
        RECT 71.000 67.900 71.900 68.200 ;
        RECT 72.900 69.200 73.300 69.900 ;
        RECT 72.900 68.800 73.800 69.200 ;
        RECT 72.900 68.200 73.300 68.800 ;
        RECT 72.900 67.900 73.800 68.200 ;
        RECT 75.000 68.000 75.400 69.900 ;
        RECT 76.600 68.000 77.000 69.900 ;
        RECT 75.000 67.900 77.000 68.000 ;
        RECT 77.400 67.900 77.800 69.900 ;
        RECT 78.200 68.500 78.600 69.500 ;
        RECT 69.400 66.100 69.800 66.200 ;
        RECT 67.000 65.800 67.800 66.100 ;
        RECT 68.600 65.800 69.800 66.100 ;
        RECT 61.400 65.700 61.700 65.800 ;
        RECT 60.700 65.400 61.700 65.700 ;
        RECT 62.600 65.600 63.000 65.800 ;
        RECT 60.700 65.100 61.000 65.400 ;
        RECT 63.900 65.100 64.200 65.800 ;
        RECT 67.400 65.600 67.800 65.800 ;
        RECT 69.400 65.100 69.700 65.800 ;
        RECT 57.100 61.100 58.100 65.100 ;
        RECT 59.800 61.400 60.200 65.100 ;
        RECT 60.600 61.700 61.000 65.100 ;
        RECT 61.400 64.800 63.400 65.100 ;
        RECT 61.400 61.400 61.800 64.800 ;
        RECT 59.800 61.100 61.800 61.400 ;
        RECT 63.000 61.100 63.400 64.800 ;
        RECT 63.800 61.100 64.200 65.100 ;
        RECT 64.600 64.800 66.600 65.100 ;
        RECT 64.600 61.100 65.000 64.800 ;
        RECT 66.200 61.100 66.600 64.800 ;
        RECT 67.000 64.800 69.000 65.100 ;
        RECT 67.000 61.100 67.400 64.800 ;
        RECT 68.600 61.100 69.000 64.800 ;
        RECT 69.400 61.100 69.800 65.100 ;
        RECT 71.000 61.100 71.400 67.900 ;
        RECT 71.800 65.100 72.200 65.200 ;
        RECT 72.600 65.100 73.000 65.200 ;
        RECT 71.800 64.800 73.000 65.100 ;
        RECT 71.800 64.400 72.200 64.800 ;
        RECT 72.600 64.400 73.000 64.800 ;
        RECT 73.400 61.100 73.800 67.900 ;
        RECT 75.100 67.700 76.900 67.900 ;
        RECT 75.400 67.200 75.800 67.400 ;
        RECT 77.400 67.200 77.700 67.900 ;
        RECT 78.200 67.400 78.500 68.500 ;
        RECT 80.300 68.000 80.700 69.500 ;
        RECT 84.300 69.200 84.700 69.900 ;
        RECT 86.700 69.200 87.100 69.900 ;
        RECT 84.300 68.800 85.000 69.200 ;
        RECT 86.700 68.800 87.400 69.200 ;
        RECT 88.600 68.900 89.000 69.900 ;
        RECT 84.300 68.200 84.700 68.800 ;
        RECT 86.700 68.200 87.100 68.800 ;
        RECT 80.300 67.700 81.100 68.000 ;
        RECT 80.700 67.500 81.100 67.700 ;
        RECT 75.000 66.900 75.800 67.200 ;
        RECT 75.000 66.800 75.400 66.900 ;
        RECT 76.500 66.800 77.800 67.200 ;
        RECT 78.200 67.100 80.300 67.400 ;
        RECT 79.800 66.900 80.300 67.100 ;
        RECT 80.800 67.200 81.100 67.500 ;
        RECT 83.800 67.900 84.700 68.200 ;
        RECT 86.200 67.900 87.100 68.200 ;
        RECT 75.000 66.100 75.400 66.200 ;
        RECT 75.800 66.100 76.200 66.600 ;
        RECT 75.000 65.800 76.200 66.100 ;
        RECT 76.500 65.100 76.800 66.800 ;
        RECT 77.400 66.100 77.800 66.200 ;
        RECT 78.200 66.100 78.600 66.600 ;
        RECT 77.400 65.800 78.600 66.100 ;
        RECT 79.800 66.500 80.500 66.900 ;
        RECT 80.800 66.800 81.800 67.200 ;
        RECT 79.800 65.500 80.100 66.500 ;
        RECT 78.200 65.200 80.100 65.500 ;
        RECT 77.400 65.100 77.800 65.200 ;
        RECT 76.300 64.800 76.800 65.100 ;
        RECT 77.100 64.800 77.800 65.100 ;
        RECT 76.300 62.200 76.700 64.800 ;
        RECT 77.100 64.200 77.400 64.800 ;
        RECT 77.000 63.800 77.400 64.200 ;
        RECT 75.800 61.800 76.700 62.200 ;
        RECT 76.300 61.100 76.700 61.800 ;
        RECT 78.200 63.500 78.500 65.200 ;
        RECT 80.800 64.900 81.100 66.800 ;
        RECT 80.300 64.600 81.100 64.900 ;
        RECT 78.200 61.500 78.600 63.500 ;
        RECT 80.300 62.200 80.700 64.600 ;
        RECT 80.300 61.800 81.000 62.200 ;
        RECT 80.300 61.100 80.700 61.800 ;
        RECT 83.800 61.100 84.200 67.900 ;
        RECT 84.600 64.400 85.000 65.200 ;
        RECT 86.200 61.100 86.600 67.900 ;
        RECT 88.700 67.200 89.000 68.900 ;
        RECT 88.600 66.800 89.000 67.200 ;
        RECT 87.000 64.400 87.400 65.200 ;
        RECT 88.700 65.100 89.000 66.800 ;
        RECT 91.000 67.100 91.400 69.900 ;
        RECT 91.800 68.000 92.200 69.900 ;
        RECT 93.400 68.000 93.800 69.900 ;
        RECT 91.800 67.900 93.800 68.000 ;
        RECT 94.200 67.900 94.600 69.900 ;
        RECT 95.800 68.800 96.200 69.900 ;
        RECT 91.900 67.700 93.700 67.900 ;
        RECT 92.200 67.200 92.600 67.400 ;
        RECT 94.200 67.200 94.500 67.900 ;
        RECT 95.900 67.200 96.200 68.800 ;
        RECT 91.800 67.100 92.600 67.200 ;
        RECT 91.000 66.900 92.600 67.100 ;
        RECT 91.000 66.800 92.200 66.900 ;
        RECT 93.300 66.800 94.600 67.200 ;
        RECT 95.800 66.800 96.200 67.200 ;
        RECT 91.000 66.100 91.400 66.800 ;
        RECT 91.800 66.100 92.200 66.200 ;
        RECT 91.000 65.800 92.200 66.100 ;
        RECT 92.600 65.800 93.000 66.600 ;
        RECT 88.600 64.700 89.500 65.100 ;
        RECT 89.100 64.100 89.500 64.700 ;
        RECT 90.200 64.800 90.600 65.200 ;
        RECT 90.200 64.100 90.500 64.800 ;
        RECT 89.100 63.800 90.500 64.100 ;
        RECT 89.100 61.100 89.500 63.800 ;
        RECT 91.000 61.100 91.400 65.800 ;
        RECT 93.300 65.100 93.600 66.800 ;
        RECT 94.200 65.100 94.600 65.200 ;
        RECT 95.900 65.100 96.200 66.800 ;
        RECT 98.200 68.900 98.600 69.900 ;
        RECT 98.200 68.200 98.500 68.900 ;
        RECT 98.200 67.800 98.600 68.200 ;
        RECT 99.000 67.800 99.400 68.600 ;
        RECT 101.400 68.000 101.800 69.900 ;
        RECT 103.000 68.000 103.400 69.900 ;
        RECT 101.400 67.900 103.400 68.000 ;
        RECT 103.800 67.900 104.200 69.900 ;
        RECT 105.900 69.200 106.300 69.900 ;
        RECT 105.400 68.800 106.300 69.200 ;
        RECT 105.900 68.200 106.300 68.800 ;
        RECT 105.400 67.900 106.300 68.200 ;
        RECT 107.000 67.900 107.400 69.900 ;
        RECT 107.800 68.000 108.200 69.900 ;
        RECT 109.400 68.000 109.800 69.900 ;
        RECT 107.800 67.900 109.800 68.000 ;
        RECT 110.200 67.900 110.600 69.900 ;
        RECT 111.000 68.000 111.400 69.900 ;
        RECT 112.600 68.000 113.000 69.900 ;
        RECT 111.000 67.900 113.000 68.000 ;
        RECT 114.200 68.800 114.600 69.900 ;
        RECT 98.200 67.200 98.500 67.800 ;
        RECT 101.500 67.700 103.300 67.900 ;
        RECT 101.800 67.200 102.200 67.400 ;
        RECT 103.800 67.200 104.100 67.900 ;
        RECT 98.200 66.800 98.600 67.200 ;
        RECT 101.400 66.900 102.200 67.200 ;
        RECT 101.400 66.800 101.800 66.900 ;
        RECT 102.900 66.800 104.200 67.200 ;
        RECT 104.600 66.800 105.000 67.600 ;
        RECT 96.600 65.400 97.000 66.200 ;
        RECT 98.200 65.100 98.500 66.800 ;
        RECT 102.200 65.800 102.600 66.600 ;
        RECT 102.900 66.100 103.200 66.800 ;
        RECT 104.600 66.100 105.000 66.200 ;
        RECT 102.900 65.800 105.000 66.100 ;
        RECT 102.900 65.100 103.200 65.800 ;
        RECT 103.800 65.100 104.200 65.200 ;
        RECT 93.100 64.800 93.600 65.100 ;
        RECT 93.900 64.800 94.600 65.100 ;
        RECT 93.100 62.200 93.500 64.800 ;
        RECT 93.900 64.200 94.200 64.800 ;
        RECT 95.800 64.700 96.700 65.100 ;
        RECT 93.800 63.800 94.200 64.200 ;
        RECT 92.600 61.800 93.500 62.200 ;
        RECT 93.100 61.100 93.500 61.800 ;
        RECT 96.300 61.100 96.700 64.700 ;
        RECT 97.700 64.700 98.600 65.100 ;
        RECT 102.700 64.800 103.200 65.100 ;
        RECT 103.500 64.800 104.200 65.100 ;
        RECT 97.700 61.100 98.100 64.700 ;
        RECT 102.700 61.100 103.100 64.800 ;
        RECT 103.500 64.200 103.800 64.800 ;
        RECT 103.400 63.800 103.800 64.200 ;
        RECT 105.400 61.100 105.800 67.900 ;
        RECT 107.100 67.200 107.400 67.900 ;
        RECT 107.900 67.700 109.700 67.900 ;
        RECT 109.000 67.200 109.400 67.400 ;
        RECT 110.300 67.200 110.600 67.900 ;
        RECT 111.100 67.700 112.900 67.900 ;
        RECT 112.200 67.200 112.600 67.400 ;
        RECT 114.200 67.200 114.500 68.800 ;
        RECT 115.000 67.800 115.400 68.600 ;
        RECT 115.800 68.000 116.200 69.900 ;
        RECT 117.400 68.000 117.800 69.900 ;
        RECT 115.800 67.900 117.800 68.000 ;
        RECT 118.200 67.900 118.600 69.900 ;
        RECT 119.800 68.900 120.200 69.900 ;
        RECT 115.900 67.700 117.700 67.900 ;
        RECT 116.200 67.200 116.600 67.400 ;
        RECT 118.200 67.200 118.500 67.900 ;
        RECT 119.000 67.800 119.400 68.600 ;
        RECT 119.900 67.200 120.200 68.900 ;
        RECT 122.700 68.200 123.100 69.900 ;
        RECT 122.200 67.900 123.100 68.200 ;
        RECT 123.800 67.900 124.200 69.900 ;
        RECT 124.600 68.000 125.000 69.900 ;
        RECT 126.200 68.000 126.600 69.900 ;
        RECT 124.600 67.900 126.600 68.000 ;
        RECT 107.000 66.800 108.300 67.200 ;
        RECT 109.000 66.900 109.800 67.200 ;
        RECT 109.400 66.800 109.800 66.900 ;
        RECT 110.200 66.800 111.500 67.200 ;
        RECT 112.200 66.900 113.000 67.200 ;
        RECT 112.600 66.800 113.000 66.900 ;
        RECT 114.200 66.800 114.600 67.200 ;
        RECT 115.000 67.100 115.400 67.200 ;
        RECT 115.800 67.100 116.600 67.200 ;
        RECT 115.000 66.900 116.600 67.100 ;
        RECT 115.000 66.800 116.200 66.900 ;
        RECT 117.300 66.800 118.600 67.200 ;
        RECT 119.800 67.100 120.200 67.200 ;
        RECT 121.400 67.100 121.800 67.600 ;
        RECT 119.800 66.800 121.800 67.100 ;
        RECT 106.200 64.400 106.600 65.200 ;
        RECT 107.000 65.100 107.400 65.200 ;
        RECT 108.000 65.100 108.300 66.800 ;
        RECT 108.600 66.100 109.000 66.600 ;
        RECT 111.200 66.100 111.500 66.800 ;
        RECT 108.600 65.800 111.500 66.100 ;
        RECT 111.800 65.800 112.200 66.600 ;
        RECT 112.600 66.100 113.000 66.200 ;
        RECT 113.400 66.100 113.800 66.200 ;
        RECT 112.600 65.800 113.800 66.100 ;
        RECT 110.200 65.100 110.600 65.200 ;
        RECT 111.200 65.100 111.500 65.800 ;
        RECT 113.400 65.400 113.800 65.800 ;
        RECT 114.200 65.100 114.500 66.800 ;
        RECT 116.600 65.800 117.000 66.600 ;
        RECT 117.300 65.100 117.600 66.800 ;
        RECT 118.200 65.100 118.600 65.200 ;
        RECT 119.900 65.100 120.200 66.800 ;
        RECT 120.600 65.400 121.000 66.200 ;
        RECT 107.000 64.800 107.700 65.100 ;
        RECT 108.000 64.800 108.500 65.100 ;
        RECT 110.200 64.800 110.900 65.100 ;
        RECT 111.200 64.800 111.700 65.100 ;
        RECT 107.400 64.200 107.700 64.800 ;
        RECT 107.400 63.800 107.800 64.200 ;
        RECT 108.100 62.200 108.500 64.800 ;
        RECT 110.600 64.200 110.900 64.800 ;
        RECT 110.600 63.800 111.000 64.200 ;
        RECT 108.100 61.800 109.000 62.200 ;
        RECT 108.100 61.100 108.500 61.800 ;
        RECT 111.300 61.100 111.700 64.800 ;
        RECT 113.700 64.700 114.600 65.100 ;
        RECT 117.100 64.800 117.600 65.100 ;
        RECT 117.900 64.800 118.600 65.100 ;
        RECT 113.700 61.100 114.100 64.700 ;
        RECT 117.100 61.100 117.500 64.800 ;
        RECT 117.900 64.200 118.200 64.800 ;
        RECT 119.800 64.700 120.700 65.100 ;
        RECT 117.800 63.800 118.200 64.200 ;
        RECT 120.300 61.100 120.700 64.700 ;
        RECT 122.200 61.100 122.600 67.900 ;
        RECT 123.900 67.200 124.200 67.900 ;
        RECT 124.700 67.700 126.500 67.900 ;
        RECT 127.000 67.800 127.400 68.600 ;
        RECT 125.800 67.200 126.200 67.400 ;
        RECT 123.800 66.800 125.100 67.200 ;
        RECT 125.800 66.900 126.600 67.200 ;
        RECT 126.200 66.800 126.600 66.900 ;
        RECT 123.000 64.400 123.400 65.200 ;
        RECT 123.800 65.100 124.200 65.200 ;
        RECT 124.800 65.100 125.100 66.800 ;
        RECT 125.400 65.800 125.800 66.600 ;
        RECT 127.000 66.100 127.400 66.200 ;
        RECT 127.800 66.100 128.200 69.900 ;
        RECT 129.900 69.200 130.300 69.900 ;
        RECT 129.900 68.800 130.600 69.200 ;
        RECT 129.900 68.200 130.300 68.800 ;
        RECT 129.400 67.900 130.300 68.200 ;
        RECT 128.600 66.800 129.000 67.600 ;
        RECT 127.000 65.800 128.200 66.100 ;
        RECT 123.800 64.800 124.500 65.100 ;
        RECT 124.800 64.800 125.300 65.100 ;
        RECT 124.200 64.200 124.500 64.800 ;
        RECT 124.200 63.800 124.600 64.200 ;
        RECT 124.900 61.100 125.300 64.800 ;
        RECT 127.800 61.100 128.200 65.800 ;
        RECT 129.400 61.100 129.800 67.900 ;
        RECT 131.000 67.800 131.400 68.600 ;
        RECT 130.200 64.400 130.600 65.200 ;
        RECT 131.800 61.100 132.200 69.900 ;
        RECT 134.100 67.900 134.900 69.900 ;
        RECT 137.900 67.900 138.700 69.900 ;
        RECT 142.400 69.200 142.800 69.900 ;
        RECT 142.400 68.800 143.400 69.200 ;
        RECT 133.400 66.400 133.800 67.200 ;
        RECT 134.300 66.200 134.600 67.900 ;
        RECT 135.000 66.800 135.400 67.200 ;
        RECT 137.400 66.800 137.800 67.200 ;
        RECT 135.000 66.600 135.300 66.800 ;
        RECT 134.900 66.200 135.300 66.600 ;
        RECT 137.500 66.600 137.800 66.800 ;
        RECT 137.500 66.200 137.900 66.600 ;
        RECT 138.200 66.200 138.500 67.900 ;
        RECT 139.000 66.400 139.400 67.200 ;
        RECT 142.400 67.100 142.800 68.800 ;
        RECT 143.800 67.900 144.200 69.900 ;
        RECT 145.400 68.900 145.800 69.900 ;
        RECT 142.400 66.900 143.300 67.100 ;
        RECT 142.500 66.800 143.300 66.900 ;
        RECT 132.600 66.100 133.000 66.200 ;
        RECT 132.600 65.800 133.400 66.100 ;
        RECT 134.200 65.800 134.600 66.200 ;
        RECT 133.000 65.600 133.400 65.800 ;
        RECT 134.300 65.700 134.600 65.800 ;
        RECT 134.300 65.400 135.300 65.700 ;
        RECT 135.800 65.400 136.200 66.200 ;
        RECT 136.600 65.400 137.000 66.200 ;
        RECT 138.200 65.800 138.600 66.200 ;
        RECT 139.800 66.100 140.200 66.200 ;
        RECT 139.400 65.800 140.200 66.100 ;
        RECT 141.400 65.800 142.200 66.200 ;
        RECT 138.200 65.700 138.500 65.800 ;
        RECT 137.500 65.400 138.500 65.700 ;
        RECT 139.400 65.600 139.800 65.800 ;
        RECT 135.000 65.100 135.300 65.400 ;
        RECT 137.500 65.200 137.800 65.400 ;
        RECT 132.600 64.800 134.600 65.100 ;
        RECT 132.600 61.100 133.000 64.800 ;
        RECT 134.200 61.400 134.600 64.800 ;
        RECT 135.000 61.700 135.400 65.100 ;
        RECT 135.800 61.400 136.200 65.100 ;
        RECT 134.200 61.100 136.200 61.400 ;
        RECT 136.600 61.400 137.000 65.100 ;
        RECT 137.400 61.700 137.800 65.200 ;
        RECT 138.200 64.800 140.200 65.100 ;
        RECT 140.600 64.800 141.000 65.600 ;
        RECT 143.000 65.200 143.300 66.800 ;
        RECT 143.800 66.200 144.100 67.900 ;
        RECT 145.400 67.800 145.700 68.900 ;
        RECT 144.500 67.500 145.700 67.800 ;
        RECT 146.200 67.800 146.600 68.600 ;
        RECT 147.100 68.200 147.500 68.600 ;
        RECT 147.000 67.800 147.400 68.200 ;
        RECT 147.800 67.900 148.200 69.900 ;
        RECT 143.800 65.800 144.200 66.200 ;
        RECT 144.500 66.000 144.800 67.500 ;
        RECT 145.300 66.800 145.800 67.200 ;
        RECT 146.200 67.100 146.500 67.800 ;
        RECT 147.900 67.100 148.200 67.900 ;
        RECT 146.200 66.800 148.200 67.100 ;
        RECT 145.200 66.400 145.600 66.800 ;
        RECT 147.000 66.100 147.400 66.200 ;
        RECT 147.900 66.100 148.200 66.800 ;
        RECT 148.600 66.400 149.000 67.200 ;
        RECT 149.400 66.100 149.800 66.200 ;
        RECT 143.000 64.800 143.400 65.200 ;
        RECT 143.800 65.100 144.100 65.800 ;
        RECT 144.500 65.700 144.900 66.000 ;
        RECT 147.000 65.800 148.200 66.100 ;
        RECT 149.000 65.800 149.800 66.100 ;
        RECT 144.500 65.600 146.600 65.700 ;
        RECT 144.600 65.400 146.600 65.600 ;
        RECT 143.800 64.800 144.500 65.100 ;
        RECT 138.200 61.400 138.600 64.800 ;
        RECT 136.600 61.100 138.600 61.400 ;
        RECT 139.800 61.100 140.200 64.800 ;
        RECT 142.200 63.800 142.600 64.600 ;
        RECT 143.000 63.500 143.300 64.800 ;
        RECT 141.500 63.200 143.300 63.500 ;
        RECT 141.500 63.100 141.800 63.200 ;
        RECT 141.400 61.100 141.800 63.100 ;
        RECT 143.000 63.100 143.300 63.200 ;
        RECT 143.000 61.100 143.400 63.100 ;
        RECT 144.100 61.100 144.500 64.800 ;
        RECT 146.200 61.100 146.600 65.400 ;
        RECT 147.100 65.100 147.400 65.800 ;
        RECT 149.000 65.600 149.400 65.800 ;
        RECT 147.000 61.100 147.400 65.100 ;
        RECT 147.800 64.800 149.800 65.100 ;
        RECT 147.800 61.100 148.200 64.800 ;
        RECT 149.400 61.100 149.800 64.800 ;
        RECT 1.400 56.100 1.800 59.900 ;
        RECT 3.000 57.900 3.400 59.900 ;
        RECT 3.100 57.800 3.400 57.900 ;
        RECT 4.600 57.900 5.000 59.900 ;
        RECT 4.600 57.800 4.900 57.900 ;
        RECT 3.100 57.500 4.900 57.800 ;
        RECT 3.800 56.400 4.200 57.200 ;
        RECT 4.600 56.200 4.900 57.500 ;
        RECT 5.700 57.200 6.100 59.900 ;
        RECT 5.400 56.800 6.100 57.200 ;
        RECT 5.700 56.200 6.100 56.800 ;
        RECT 2.200 56.100 2.600 56.200 ;
        RECT 1.400 55.800 2.600 56.100 ;
        RECT 0.600 52.400 1.000 53.200 ;
        RECT 1.400 51.100 1.800 55.800 ;
        RECT 2.200 55.400 2.600 55.800 ;
        RECT 4.600 55.800 5.000 56.200 ;
        RECT 5.400 55.900 6.100 56.200 ;
        RECT 3.000 54.800 3.800 55.200 ;
        RECT 4.600 54.200 4.900 55.800 ;
        RECT 4.100 54.100 4.900 54.200 ;
        RECT 4.000 53.900 4.900 54.100 ;
        RECT 5.400 55.200 5.700 55.900 ;
        RECT 7.800 55.600 8.200 59.900 ;
        RECT 8.600 56.800 9.400 57.200 ;
        RECT 9.000 56.200 9.300 56.800 ;
        RECT 9.700 56.200 10.100 59.900 ;
        RECT 12.900 59.200 13.300 59.900 ;
        RECT 12.900 58.800 13.800 59.200 ;
        RECT 11.800 56.800 12.600 57.200 ;
        RECT 12.200 56.200 12.500 56.800 ;
        RECT 12.900 56.200 13.300 58.800 ;
        RECT 8.600 55.900 9.300 56.200 ;
        RECT 9.600 55.900 10.100 56.200 ;
        RECT 11.800 55.900 12.500 56.200 ;
        RECT 12.800 55.900 13.300 56.200 ;
        RECT 15.000 56.200 15.400 59.900 ;
        RECT 16.600 56.200 17.000 59.900 ;
        RECT 15.000 55.900 17.000 56.200 ;
        RECT 17.400 55.900 17.800 59.900 ;
        RECT 19.000 57.900 19.400 59.900 ;
        RECT 19.100 57.800 19.400 57.900 ;
        RECT 20.600 57.900 21.000 59.900 ;
        RECT 21.400 57.900 21.800 59.900 ;
        RECT 20.600 57.800 20.900 57.900 ;
        RECT 19.100 57.500 20.900 57.800 ;
        RECT 19.800 56.400 20.200 57.200 ;
        RECT 20.600 56.200 20.900 57.500 ;
        RECT 21.500 57.800 21.800 57.900 ;
        RECT 23.000 57.900 23.400 59.900 ;
        RECT 23.000 57.800 23.300 57.900 ;
        RECT 24.600 57.800 25.000 59.900 ;
        RECT 26.200 57.900 26.600 59.900 ;
        RECT 26.200 57.800 26.500 57.900 ;
        RECT 21.500 57.500 23.300 57.800 ;
        RECT 24.700 57.500 26.500 57.800 ;
        RECT 21.500 56.200 21.800 57.500 ;
        RECT 22.200 56.400 22.600 57.200 ;
        RECT 24.700 56.200 25.000 57.500 ;
        RECT 25.400 56.400 25.800 57.200 ;
        RECT 8.600 55.800 9.000 55.900 ;
        RECT 6.200 55.400 8.200 55.600 ;
        RECT 6.100 55.300 8.200 55.400 ;
        RECT 5.400 54.800 5.800 55.200 ;
        RECT 6.100 55.000 6.500 55.300 ;
        RECT 4.000 52.200 4.400 53.900 ;
        RECT 3.800 51.800 4.400 52.200 ;
        RECT 4.000 51.100 4.400 51.800 ;
        RECT 5.400 53.100 5.700 54.800 ;
        RECT 6.100 53.500 6.400 55.000 ;
        RECT 6.800 54.200 7.200 54.600 ;
        RECT 9.600 54.200 9.900 55.900 ;
        RECT 11.800 55.800 12.200 55.900 ;
        RECT 10.200 55.100 10.600 55.200 ;
        RECT 11.800 55.100 12.100 55.800 ;
        RECT 10.200 54.800 12.100 55.100 ;
        RECT 10.200 54.400 10.600 54.800 ;
        RECT 12.800 54.200 13.100 55.900 ;
        RECT 15.400 55.200 15.800 55.400 ;
        RECT 17.400 55.200 17.700 55.900 ;
        RECT 18.200 55.400 18.600 56.200 ;
        RECT 20.600 55.800 21.000 56.200 ;
        RECT 21.400 55.800 21.800 56.200 ;
        RECT 13.400 54.400 13.800 55.200 ;
        RECT 15.000 54.900 15.800 55.200 ;
        RECT 16.600 54.900 17.800 55.200 ;
        RECT 15.000 54.800 15.400 54.900 ;
        RECT 6.900 53.800 7.400 54.200 ;
        RECT 8.600 53.800 9.900 54.200 ;
        RECT 11.000 54.100 11.400 54.200 ;
        RECT 10.600 53.800 11.400 54.100 ;
        RECT 11.800 53.800 13.100 54.200 ;
        RECT 14.200 54.100 14.600 54.200 ;
        RECT 13.800 53.800 14.600 54.100 ;
        RECT 15.800 53.800 16.200 54.600 ;
        RECT 6.100 53.200 7.300 53.500 ;
        RECT 5.400 51.100 5.800 53.100 ;
        RECT 7.000 52.100 7.300 53.200 ;
        RECT 7.800 52.400 8.200 53.200 ;
        RECT 8.700 53.100 9.000 53.800 ;
        RECT 10.600 53.600 11.000 53.800 ;
        RECT 9.500 53.100 11.300 53.300 ;
        RECT 11.900 53.100 12.200 53.800 ;
        RECT 13.800 53.600 14.200 53.800 ;
        RECT 12.700 53.100 14.500 53.300 ;
        RECT 16.600 53.100 16.900 54.900 ;
        RECT 17.400 54.800 17.800 54.900 ;
        RECT 19.000 54.800 19.800 55.200 ;
        RECT 20.600 54.200 20.900 55.800 ;
        RECT 20.100 54.100 20.900 54.200 ;
        RECT 20.000 53.900 20.900 54.100 ;
        RECT 21.500 54.200 21.800 55.800 ;
        RECT 23.800 55.400 24.200 56.200 ;
        RECT 24.600 55.800 25.000 56.200 ;
        RECT 22.600 54.800 23.400 55.200 ;
        RECT 24.700 54.200 25.000 55.800 ;
        RECT 27.000 55.400 27.400 56.200 ;
        RECT 27.800 55.900 28.200 59.900 ;
        RECT 28.600 56.200 29.000 59.900 ;
        RECT 30.200 56.200 30.600 59.900 ;
        RECT 31.800 57.800 32.200 59.900 ;
        RECT 33.400 57.900 33.800 59.900 ;
        RECT 35.000 57.900 35.400 59.900 ;
        RECT 33.400 57.800 33.700 57.900 ;
        RECT 31.900 57.500 33.700 57.800 ;
        RECT 35.100 57.800 35.400 57.900 ;
        RECT 36.600 57.900 37.000 59.900 ;
        RECT 36.600 57.800 36.900 57.900 ;
        RECT 35.100 57.500 36.900 57.800 ;
        RECT 32.600 56.400 33.000 57.200 ;
        RECT 33.400 56.200 33.700 57.500 ;
        RECT 35.800 56.400 36.200 57.200 ;
        RECT 36.600 56.200 36.900 57.500 ;
        RECT 28.600 55.900 30.600 56.200 ;
        RECT 27.900 55.200 28.200 55.900 ;
        RECT 31.000 55.400 31.400 56.200 ;
        RECT 33.400 55.800 33.800 56.200 ;
        RECT 29.800 55.200 30.200 55.400 ;
        RECT 25.800 54.800 26.600 55.200 ;
        RECT 27.800 54.900 29.000 55.200 ;
        RECT 29.800 54.900 30.600 55.200 ;
        RECT 27.800 54.800 28.200 54.900 ;
        RECT 21.500 54.100 22.300 54.200 ;
        RECT 24.700 54.100 25.500 54.200 ;
        RECT 21.500 53.900 22.400 54.100 ;
        RECT 24.700 53.900 25.600 54.100 ;
        RECT 7.000 51.100 7.400 52.100 ;
        RECT 8.600 51.100 9.000 53.100 ;
        RECT 9.400 53.000 11.400 53.100 ;
        RECT 9.400 51.100 9.800 53.000 ;
        RECT 11.000 51.100 11.400 53.000 ;
        RECT 11.800 51.100 12.200 53.100 ;
        RECT 12.600 53.000 14.600 53.100 ;
        RECT 12.600 51.100 13.000 53.000 ;
        RECT 14.200 51.100 14.600 53.000 ;
        RECT 16.600 51.100 17.000 53.100 ;
        RECT 17.400 52.800 17.800 53.200 ;
        RECT 17.300 52.400 17.700 52.800 ;
        RECT 20.000 51.100 20.400 53.900 ;
        RECT 22.000 51.100 22.400 53.900 ;
        RECT 25.200 51.100 25.600 53.900 ;
        RECT 27.800 52.800 28.200 53.200 ;
        RECT 28.700 53.100 29.000 54.900 ;
        RECT 30.200 54.800 30.600 54.900 ;
        RECT 31.800 54.800 32.600 55.200 ;
        RECT 29.400 53.800 29.800 54.600 ;
        RECT 33.400 54.200 33.700 55.800 ;
        RECT 34.200 55.400 34.600 56.200 ;
        RECT 36.600 55.800 37.000 56.200 ;
        RECT 38.700 55.900 39.700 59.900 ;
        RECT 41.400 59.600 43.400 59.900 ;
        RECT 41.400 55.900 41.800 59.600 ;
        RECT 42.200 55.900 42.600 59.300 ;
        RECT 43.000 56.200 43.400 59.600 ;
        RECT 44.600 56.200 45.000 59.900 ;
        RECT 43.000 55.900 45.000 56.200 ;
        RECT 45.400 55.900 45.800 59.900 ;
        RECT 46.200 56.200 46.600 59.900 ;
        RECT 47.800 56.200 48.200 59.900 ;
        RECT 49.400 59.100 49.800 59.200 ;
        RECT 50.200 59.100 50.600 59.900 ;
        RECT 49.400 58.800 50.600 59.100 ;
        RECT 46.200 55.900 48.200 56.200 ;
        RECT 35.000 54.800 35.800 55.200 ;
        RECT 36.600 54.200 36.900 55.800 ;
        RECT 38.200 54.400 38.600 55.200 ;
        RECT 39.000 54.200 39.300 55.900 ;
        RECT 42.300 55.600 42.600 55.900 ;
        RECT 39.800 54.400 40.200 55.200 ;
        RECT 41.400 54.800 41.800 55.600 ;
        RECT 42.300 55.300 43.300 55.600 ;
        RECT 43.000 55.200 43.300 55.300 ;
        RECT 44.200 55.200 44.600 55.400 ;
        RECT 45.500 55.200 45.800 55.900 ;
        RECT 47.400 55.200 47.800 55.400 ;
        RECT 43.000 54.800 43.400 55.200 ;
        RECT 44.200 54.900 45.000 55.200 ;
        RECT 44.600 54.800 45.000 54.900 ;
        RECT 45.400 54.900 46.600 55.200 ;
        RECT 47.400 55.100 48.200 55.200 ;
        RECT 50.200 55.100 50.600 58.800 ;
        RECT 51.800 55.900 52.200 59.900 ;
        RECT 52.600 56.200 53.000 59.900 ;
        RECT 54.200 56.200 54.600 59.900 ;
        RECT 56.300 59.200 56.700 59.900 ;
        RECT 55.800 58.800 56.700 59.200 ;
        RECT 56.300 56.300 56.700 58.800 ;
        RECT 52.600 55.900 54.600 56.200 ;
        RECT 55.800 55.900 56.700 56.300 ;
        RECT 57.400 55.900 57.800 59.900 ;
        RECT 58.200 56.200 58.600 59.900 ;
        RECT 59.800 56.200 60.200 59.900 ;
        RECT 58.200 55.900 60.200 56.200 ;
        RECT 51.900 55.200 52.200 55.900 ;
        RECT 53.800 55.200 54.200 55.400 ;
        RECT 47.400 54.900 50.600 55.100 ;
        RECT 45.400 54.800 45.800 54.900 ;
        RECT 32.900 54.100 33.700 54.200 ;
        RECT 36.100 54.100 36.900 54.200 ;
        RECT 32.800 53.900 33.700 54.100 ;
        RECT 36.000 53.900 36.900 54.100 ;
        RECT 37.400 54.100 37.800 54.200 ;
        RECT 39.000 54.100 39.400 54.200 ;
        RECT 40.600 54.100 41.000 54.600 ;
        RECT 41.400 54.100 41.800 54.200 ;
        RECT 27.900 52.400 28.300 52.800 ;
        RECT 28.600 51.100 29.000 53.100 ;
        RECT 32.800 51.100 33.200 53.900 ;
        RECT 36.000 51.100 36.400 53.900 ;
        RECT 37.400 53.800 38.200 54.100 ;
        RECT 39.000 53.800 40.200 54.100 ;
        RECT 40.600 53.800 41.800 54.100 ;
        RECT 37.800 53.600 38.200 53.800 ;
        RECT 37.500 53.100 39.300 53.300 ;
        RECT 39.900 53.100 40.200 53.800 ;
        RECT 43.000 53.200 43.300 54.800 ;
        RECT 46.300 53.200 46.600 54.900 ;
        RECT 47.800 54.800 50.600 54.900 ;
        RECT 51.000 55.100 51.400 55.200 ;
        RECT 51.800 55.100 53.000 55.200 ;
        RECT 51.000 54.900 53.000 55.100 ;
        RECT 53.800 54.900 54.600 55.200 ;
        RECT 51.000 54.800 52.200 54.900 ;
        RECT 47.000 53.800 47.400 54.600 ;
        RECT 42.200 53.100 43.300 53.200 ;
        RECT 37.400 53.000 39.400 53.100 ;
        RECT 37.400 51.100 37.800 53.000 ;
        RECT 39.000 51.400 39.400 53.000 ;
        RECT 39.800 51.700 40.200 53.100 ;
        RECT 40.600 51.400 41.000 53.100 ;
        RECT 42.200 52.800 43.500 53.100 ;
        RECT 45.400 52.800 45.800 53.200 ;
        RECT 39.000 51.100 41.000 51.400 ;
        RECT 42.700 51.100 43.500 52.800 ;
        RECT 45.500 52.400 45.900 52.800 ;
        RECT 46.200 51.100 46.600 53.200 ;
        RECT 50.200 51.100 50.600 54.800 ;
        RECT 51.000 53.400 51.400 54.200 ;
        RECT 51.800 52.800 52.200 53.200 ;
        RECT 52.700 53.100 53.000 54.900 ;
        RECT 54.200 54.800 54.600 54.900 ;
        RECT 55.900 54.200 56.200 55.900 ;
        RECT 56.600 54.800 57.000 55.600 ;
        RECT 57.500 55.200 57.800 55.900 ;
        RECT 59.400 55.200 59.800 55.400 ;
        RECT 57.400 54.900 58.600 55.200 ;
        RECT 59.400 54.900 60.200 55.200 ;
        RECT 57.400 54.800 57.800 54.900 ;
        RECT 55.800 53.800 56.200 54.200 ;
        RECT 51.900 52.400 52.300 52.800 ;
        RECT 52.600 51.100 53.000 53.100 ;
        RECT 55.000 52.400 55.400 53.200 ;
        RECT 55.900 52.100 56.200 53.800 ;
        RECT 57.400 52.800 57.800 53.200 ;
        RECT 58.300 53.100 58.600 54.900 ;
        RECT 59.800 54.800 60.200 54.900 ;
        RECT 60.600 53.400 61.000 54.200 ;
        RECT 57.500 52.400 57.900 52.800 ;
        RECT 55.800 51.100 56.200 52.100 ;
        RECT 58.200 51.100 58.600 53.100 ;
        RECT 61.400 53.100 61.800 59.900 ;
        RECT 63.800 55.600 64.200 59.900 ;
        RECT 65.400 55.600 65.800 59.900 ;
        RECT 68.300 56.300 68.700 59.900 ;
        RECT 70.700 56.300 71.100 59.900 ;
        RECT 67.800 55.900 68.700 56.300 ;
        RECT 70.200 55.900 71.100 56.300 ;
        RECT 63.800 55.200 65.800 55.600 ;
        RECT 63.000 53.400 63.400 54.200 ;
        RECT 65.400 53.800 65.800 55.200 ;
        RECT 67.900 54.200 68.200 55.900 ;
        RECT 68.600 54.800 69.000 55.600 ;
        RECT 70.300 54.200 70.600 55.900 ;
        RECT 71.000 55.100 71.400 55.600 ;
        RECT 71.800 55.100 72.200 59.900 ;
        RECT 73.700 56.300 74.100 59.900 ;
        RECT 73.700 55.900 74.600 56.300 ;
        RECT 71.000 54.800 72.200 55.100 ;
        RECT 73.400 54.800 73.800 55.600 ;
        RECT 67.800 53.800 68.200 54.200 ;
        RECT 70.200 54.100 70.600 54.200 ;
        RECT 70.200 53.800 71.300 54.100 ;
        RECT 63.800 53.400 65.800 53.800 ;
        RECT 61.400 52.800 62.300 53.100 ;
        RECT 61.900 51.100 62.300 52.800 ;
        RECT 63.800 51.100 64.200 53.400 ;
        RECT 65.400 51.100 65.800 53.400 ;
        RECT 67.000 52.400 67.400 53.200 ;
        RECT 67.900 52.200 68.200 53.800 ;
        RECT 69.400 52.400 69.800 53.200 ;
        RECT 67.800 51.100 68.200 52.200 ;
        RECT 70.300 52.100 70.600 53.800 ;
        RECT 71.000 53.200 71.300 53.800 ;
        RECT 71.000 52.800 71.400 53.200 ;
        RECT 70.200 51.100 70.600 52.100 ;
        RECT 71.800 51.100 72.200 54.800 ;
        RECT 74.200 54.200 74.500 55.900 ;
        RECT 74.200 53.800 74.600 54.200 ;
        RECT 72.600 53.100 73.000 53.200 ;
        RECT 74.200 53.100 74.500 53.800 ;
        RECT 72.600 52.800 74.500 53.100 ;
        RECT 72.600 52.400 73.000 52.800 ;
        RECT 74.200 52.100 74.500 52.800 ;
        RECT 75.000 52.400 75.400 53.200 ;
        RECT 74.200 51.100 74.600 52.100 ;
        RECT 75.800 51.100 76.200 59.900 ;
        RECT 78.500 57.200 78.900 59.900 ;
        RECT 77.800 56.800 78.200 57.200 ;
        RECT 78.500 56.800 79.400 57.200 ;
        RECT 77.800 56.200 78.100 56.800 ;
        RECT 78.500 56.200 78.900 56.800 ;
        RECT 77.400 55.900 78.100 56.200 ;
        RECT 78.400 55.900 78.900 56.200 ;
        RECT 80.600 56.100 81.000 56.200 ;
        RECT 81.400 56.100 81.800 59.900 ;
        RECT 77.400 55.800 77.800 55.900 ;
        RECT 78.400 54.200 78.700 55.900 ;
        RECT 80.600 55.800 81.800 56.100 ;
        RECT 83.300 56.300 83.700 59.900 ;
        RECT 83.300 55.900 84.200 56.300 ;
        RECT 86.700 56.200 87.100 59.900 ;
        RECT 87.400 56.800 87.800 57.200 ;
        RECT 87.500 56.200 87.800 56.800 ;
        RECT 86.700 55.900 87.200 56.200 ;
        RECT 87.500 55.900 88.200 56.200 ;
        RECT 79.000 55.100 79.400 55.200 ;
        RECT 79.000 54.800 80.900 55.100 ;
        RECT 79.000 54.400 79.400 54.800 ;
        RECT 80.600 54.200 80.900 54.800 ;
        RECT 77.400 53.800 78.700 54.200 ;
        RECT 79.800 54.100 80.200 54.200 ;
        RECT 79.400 53.800 80.200 54.100 ;
        RECT 77.500 53.100 77.800 53.800 ;
        RECT 79.400 53.600 79.800 53.800 ;
        RECT 80.600 53.400 81.000 54.200 ;
        RECT 78.300 53.100 80.100 53.300 ;
        RECT 81.400 53.100 81.800 55.800 ;
        RECT 83.000 54.800 83.400 55.600 ;
        RECT 83.800 54.200 84.100 55.900 ;
        RECT 86.200 54.400 86.600 55.200 ;
        RECT 86.900 54.200 87.200 55.900 ;
        RECT 87.800 55.800 88.200 55.900 ;
        RECT 88.600 54.800 89.000 55.200 ;
        RECT 83.800 53.800 84.200 54.200 ;
        RECT 85.400 54.100 85.800 54.200 ;
        RECT 86.900 54.100 88.200 54.200 ;
        RECT 88.600 54.100 88.900 54.800 ;
        RECT 85.400 53.800 86.200 54.100 ;
        RECT 86.900 53.800 88.900 54.100 ;
        RECT 77.400 51.100 77.800 53.100 ;
        RECT 78.200 53.000 80.200 53.100 ;
        RECT 78.200 51.100 78.600 53.000 ;
        RECT 79.800 51.100 80.200 53.000 ;
        RECT 81.400 52.800 82.300 53.100 ;
        RECT 81.900 51.100 82.300 52.800 ;
        RECT 83.800 52.200 84.100 53.800 ;
        RECT 85.800 53.600 86.200 53.800 ;
        RECT 85.500 53.100 87.300 53.300 ;
        RECT 87.800 53.100 88.100 53.800 ;
        RECT 88.600 53.100 89.000 53.200 ;
        RECT 85.400 53.000 87.400 53.100 ;
        RECT 83.800 51.100 84.200 52.200 ;
        RECT 85.400 51.100 85.800 53.000 ;
        RECT 87.000 51.100 87.400 53.000 ;
        RECT 87.800 52.800 89.000 53.100 ;
        RECT 87.800 51.100 88.200 52.800 ;
        RECT 88.600 52.400 89.000 52.800 ;
        RECT 89.400 51.100 89.800 59.900 ;
        RECT 91.500 56.200 91.900 59.900 ;
        RECT 92.200 56.800 92.600 57.200 ;
        RECT 92.300 56.200 92.600 56.800 ;
        RECT 94.700 56.200 95.100 59.900 ;
        RECT 95.400 56.800 95.800 57.200 ;
        RECT 95.500 56.200 95.800 56.800 ;
        RECT 97.900 56.300 98.300 59.900 ;
        RECT 91.500 55.900 92.000 56.200 ;
        RECT 92.300 55.900 93.000 56.200 ;
        RECT 94.700 55.900 95.200 56.200 ;
        RECT 95.500 55.900 96.200 56.200 ;
        RECT 97.400 55.900 98.300 56.300 ;
        RECT 101.900 56.200 102.300 59.900 ;
        RECT 102.600 56.800 103.000 57.200 ;
        RECT 102.700 56.200 103.000 56.800 ;
        RECT 91.000 54.400 91.400 55.200 ;
        RECT 91.700 54.200 92.000 55.900 ;
        RECT 92.600 55.800 93.000 55.900 ;
        RECT 94.200 54.400 94.600 55.200 ;
        RECT 94.900 54.200 95.200 55.900 ;
        RECT 95.800 55.800 96.200 55.900 ;
        RECT 96.600 55.100 97.000 55.200 ;
        RECT 97.500 55.100 97.800 55.900 ;
        RECT 101.400 55.800 102.400 56.200 ;
        RECT 102.700 56.100 103.400 56.200 ;
        RECT 104.600 56.100 105.000 59.900 ;
        RECT 106.700 56.300 107.100 59.900 ;
        RECT 102.700 55.900 105.000 56.100 ;
        RECT 106.200 55.900 107.100 56.300 ;
        RECT 107.800 55.900 108.200 59.900 ;
        RECT 108.600 56.200 109.000 59.900 ;
        RECT 110.200 56.200 110.600 59.900 ;
        RECT 108.600 55.900 110.600 56.200 ;
        RECT 112.300 56.200 112.700 59.900 ;
        RECT 113.000 56.800 113.400 57.200 ;
        RECT 113.100 56.200 113.400 56.800 ;
        RECT 112.300 55.900 112.800 56.200 ;
        RECT 113.100 55.900 113.800 56.200 ;
        RECT 103.000 55.800 105.000 55.900 ;
        RECT 96.600 54.800 97.800 55.100 ;
        RECT 98.200 54.800 98.600 55.600 ;
        RECT 97.500 54.200 97.800 54.800 ;
        RECT 101.400 54.400 101.800 55.200 ;
        RECT 102.100 54.200 102.400 55.800 ;
        RECT 90.200 54.100 90.600 54.200 ;
        RECT 90.200 53.800 91.000 54.100 ;
        RECT 91.700 53.800 93.000 54.200 ;
        RECT 93.400 54.100 93.800 54.200 ;
        RECT 93.400 53.800 94.200 54.100 ;
        RECT 94.900 53.800 96.200 54.200 ;
        RECT 97.400 53.800 97.800 54.200 ;
        RECT 100.600 54.100 101.000 54.200 ;
        RECT 100.600 53.800 101.400 54.100 ;
        RECT 102.100 53.800 103.400 54.200 ;
        RECT 104.600 54.100 105.000 55.800 ;
        RECT 105.400 55.100 105.800 55.200 ;
        RECT 106.300 55.100 106.600 55.900 ;
        RECT 105.400 54.800 106.600 55.100 ;
        RECT 107.000 54.800 107.400 55.600 ;
        RECT 107.900 55.200 108.200 55.900 ;
        RECT 109.800 55.200 110.200 55.400 ;
        RECT 107.800 54.900 109.000 55.200 ;
        RECT 109.800 54.900 110.600 55.200 ;
        RECT 107.800 54.800 108.200 54.900 ;
        RECT 106.300 54.200 106.600 54.800 ;
        RECT 105.400 54.100 105.800 54.200 ;
        RECT 104.600 53.800 105.800 54.100 ;
        RECT 106.200 53.800 106.600 54.200 ;
        RECT 90.600 53.600 91.000 53.800 ;
        RECT 90.300 53.100 92.100 53.300 ;
        RECT 92.600 53.100 92.900 53.800 ;
        RECT 93.800 53.600 94.200 53.800 ;
        RECT 93.500 53.100 95.300 53.300 ;
        RECT 95.800 53.100 96.100 53.800 ;
        RECT 96.600 53.100 97.000 53.200 ;
        RECT 90.200 53.000 92.200 53.100 ;
        RECT 90.200 51.100 90.600 53.000 ;
        RECT 91.800 51.100 92.200 53.000 ;
        RECT 92.600 51.100 93.000 53.100 ;
        RECT 93.400 53.000 95.400 53.100 ;
        RECT 93.400 51.100 93.800 53.000 ;
        RECT 95.000 51.100 95.400 53.000 ;
        RECT 95.800 52.800 97.000 53.100 ;
        RECT 95.800 51.100 96.200 52.800 ;
        RECT 96.600 52.400 97.000 52.800 ;
        RECT 97.500 52.100 97.800 53.800 ;
        RECT 101.000 53.600 101.400 53.800 ;
        RECT 100.700 53.100 102.500 53.300 ;
        RECT 103.000 53.100 103.300 53.800 ;
        RECT 97.400 51.100 97.800 52.100 ;
        RECT 100.600 53.000 102.600 53.100 ;
        RECT 100.600 51.100 101.000 53.000 ;
        RECT 102.200 51.100 102.600 53.000 ;
        RECT 103.000 51.100 103.400 53.100 ;
        RECT 103.800 52.400 104.200 53.200 ;
        RECT 104.600 51.100 105.000 53.800 ;
        RECT 105.400 52.400 105.800 53.200 ;
        RECT 106.300 52.100 106.600 53.800 ;
        RECT 107.800 52.800 108.200 53.200 ;
        RECT 108.700 53.100 109.000 54.900 ;
        RECT 110.200 54.800 110.600 54.900 ;
        RECT 109.400 53.800 109.800 54.600 ;
        RECT 111.800 54.400 112.200 55.200 ;
        RECT 112.500 54.200 112.800 55.900 ;
        RECT 113.400 55.800 113.800 55.900 ;
        RECT 111.000 54.100 111.400 54.200 ;
        RECT 111.000 53.800 111.800 54.100 ;
        RECT 112.500 53.800 113.800 54.200 ;
        RECT 111.400 53.600 111.800 53.800 ;
        RECT 111.100 53.100 112.900 53.300 ;
        RECT 113.400 53.100 113.700 53.800 ;
        RECT 114.200 53.100 114.600 53.200 ;
        RECT 107.900 52.400 108.300 52.800 ;
        RECT 106.200 51.100 106.600 52.100 ;
        RECT 108.600 51.100 109.000 53.100 ;
        RECT 111.000 53.000 113.000 53.100 ;
        RECT 111.000 51.100 111.400 53.000 ;
        RECT 112.600 51.100 113.000 53.000 ;
        RECT 113.400 52.800 114.600 53.100 ;
        RECT 113.400 51.100 113.800 52.800 ;
        RECT 114.200 52.400 114.600 52.800 ;
        RECT 115.000 51.100 115.400 59.900 ;
        RECT 117.100 59.200 117.500 59.900 ;
        RECT 116.600 58.800 117.500 59.200 ;
        RECT 117.100 56.200 117.500 58.800 ;
        RECT 117.800 56.800 118.200 57.200 ;
        RECT 117.900 56.200 118.200 56.800 ;
        RECT 117.100 55.900 117.600 56.200 ;
        RECT 117.900 55.900 118.600 56.200 ;
        RECT 116.600 54.400 117.000 55.200 ;
        RECT 117.300 54.200 117.600 55.900 ;
        RECT 118.200 55.800 118.600 55.900 ;
        RECT 115.800 54.100 116.200 54.200 ;
        RECT 115.800 53.800 116.600 54.100 ;
        RECT 117.300 53.800 118.600 54.200 ;
        RECT 116.200 53.600 116.600 53.800 ;
        RECT 115.900 53.100 117.700 53.300 ;
        RECT 118.200 53.100 118.500 53.800 ;
        RECT 119.000 53.400 119.400 54.200 ;
        RECT 119.800 53.100 120.200 59.900 ;
        RECT 120.600 55.800 121.000 56.600 ;
        RECT 121.700 56.300 122.100 59.900 ;
        RECT 121.700 55.900 122.600 56.300 ;
        RECT 123.800 56.200 124.200 59.900 ;
        RECT 125.400 56.200 125.800 59.900 ;
        RECT 123.800 55.900 125.800 56.200 ;
        RECT 126.200 55.900 126.600 59.900 ;
        RECT 128.300 56.200 128.700 59.900 ;
        RECT 128.300 55.900 128.800 56.200 ;
        RECT 130.200 55.900 130.600 59.900 ;
        RECT 131.000 56.200 131.400 59.900 ;
        RECT 132.600 56.200 133.000 59.900 ;
        RECT 134.200 57.900 134.600 59.900 ;
        RECT 134.300 57.800 134.600 57.900 ;
        RECT 135.800 57.900 136.200 59.900 ;
        RECT 135.800 57.800 136.100 57.900 ;
        RECT 134.300 57.500 136.100 57.800 ;
        RECT 135.000 56.400 135.400 57.200 ;
        RECT 135.800 56.200 136.100 57.500 ;
        RECT 131.000 55.900 133.000 56.200 ;
        RECT 122.200 55.800 122.600 55.900 ;
        RECT 121.400 54.800 121.800 55.600 ;
        RECT 122.200 54.200 122.500 55.800 ;
        RECT 124.200 55.200 124.600 55.400 ;
        RECT 126.200 55.200 126.500 55.900 ;
        RECT 123.800 54.900 124.600 55.200 ;
        RECT 125.400 54.900 126.600 55.200 ;
        RECT 123.800 54.800 124.200 54.900 ;
        RECT 122.200 53.800 122.600 54.200 ;
        RECT 124.600 53.800 125.000 54.600 ;
        RECT 115.800 53.000 117.800 53.100 ;
        RECT 115.800 51.100 116.200 53.000 ;
        RECT 117.400 51.100 117.800 53.000 ;
        RECT 118.200 51.100 118.600 53.100 ;
        RECT 119.800 52.800 120.700 53.100 ;
        RECT 120.300 52.200 120.700 52.800 ;
        RECT 119.800 51.800 120.700 52.200 ;
        RECT 120.300 51.100 120.700 51.800 ;
        RECT 122.200 52.100 122.500 53.800 ;
        RECT 125.400 53.200 125.700 54.900 ;
        RECT 126.200 54.800 126.600 54.900 ;
        RECT 127.800 54.400 128.200 55.200 ;
        RECT 128.500 54.200 128.800 55.900 ;
        RECT 130.300 55.200 130.600 55.900 ;
        RECT 133.400 55.400 133.800 56.200 ;
        RECT 135.800 55.800 136.200 56.200 ;
        RECT 132.200 55.200 132.600 55.400 ;
        RECT 130.200 54.900 131.400 55.200 ;
        RECT 132.200 54.900 133.000 55.200 ;
        RECT 130.200 54.800 130.600 54.900 ;
        RECT 127.000 54.100 127.400 54.200 ;
        RECT 127.000 53.800 127.800 54.100 ;
        RECT 128.500 53.800 129.800 54.200 ;
        RECT 127.400 53.600 127.800 53.800 ;
        RECT 123.000 52.400 123.400 53.200 ;
        RECT 122.200 51.100 122.600 52.100 ;
        RECT 125.400 51.100 125.800 53.200 ;
        RECT 126.200 52.800 126.600 53.200 ;
        RECT 127.100 53.100 128.900 53.300 ;
        RECT 129.400 53.100 129.700 53.800 ;
        RECT 130.200 53.100 130.600 53.200 ;
        RECT 131.100 53.100 131.400 54.900 ;
        RECT 132.600 54.800 133.000 54.900 ;
        RECT 134.200 54.800 135.000 55.200 ;
        RECT 131.800 53.800 132.200 54.600 ;
        RECT 135.800 54.200 136.100 55.800 ;
        RECT 135.300 54.100 136.100 54.200 ;
        RECT 135.200 53.900 136.100 54.100 ;
        RECT 127.000 53.000 129.000 53.100 ;
        RECT 126.100 52.400 126.500 52.800 ;
        RECT 127.000 51.100 127.400 53.000 ;
        RECT 128.600 51.100 129.000 53.000 ;
        RECT 129.400 52.800 130.600 53.100 ;
        RECT 129.400 51.100 129.800 52.800 ;
        RECT 130.300 52.400 130.700 52.800 ;
        RECT 131.000 51.100 131.400 53.100 ;
        RECT 135.200 51.100 135.600 53.900 ;
        RECT 136.600 53.400 137.000 54.200 ;
        RECT 137.400 51.100 137.800 59.900 ;
        RECT 140.300 56.200 140.700 59.900 ;
        RECT 141.000 56.800 141.400 57.200 ;
        RECT 141.100 56.200 141.400 56.800 ;
        RECT 143.500 56.300 143.900 59.900 ;
        RECT 144.900 59.200 145.300 59.900 ;
        RECT 144.600 58.800 145.300 59.200 ;
        RECT 140.300 55.900 140.800 56.200 ;
        RECT 141.100 55.900 141.800 56.200 ;
        RECT 143.000 55.900 143.900 56.300 ;
        RECT 144.900 56.300 145.300 58.800 ;
        RECT 144.900 55.900 145.800 56.300 ;
        RECT 139.000 55.100 139.400 55.200 ;
        RECT 139.800 55.100 140.200 55.200 ;
        RECT 139.000 54.800 140.200 55.100 ;
        RECT 139.800 54.400 140.200 54.800 ;
        RECT 140.500 54.200 140.800 55.900 ;
        RECT 141.400 55.800 141.800 55.900 ;
        RECT 141.400 55.100 141.700 55.800 ;
        RECT 143.100 55.100 143.400 55.900 ;
        RECT 141.400 54.800 143.400 55.100 ;
        RECT 143.800 55.100 144.200 55.600 ;
        RECT 144.600 55.100 145.000 55.600 ;
        RECT 143.800 54.800 145.000 55.100 ;
        RECT 143.100 54.200 143.400 54.800 ;
        RECT 140.500 53.800 141.800 54.200 ;
        RECT 142.200 54.100 142.600 54.200 ;
        RECT 143.000 54.100 143.400 54.200 ;
        RECT 142.200 53.800 143.400 54.100 ;
        RECT 139.100 53.100 140.900 53.300 ;
        RECT 141.400 53.100 141.700 53.800 ;
        RECT 139.000 53.000 141.000 53.100 ;
        RECT 139.000 51.100 139.400 53.000 ;
        RECT 140.600 51.100 141.000 53.000 ;
        RECT 141.400 51.100 141.800 53.100 ;
        RECT 142.200 52.400 142.600 53.200 ;
        RECT 143.100 52.100 143.400 53.800 ;
        RECT 143.000 51.100 143.400 52.100 ;
        RECT 145.400 54.200 145.700 55.900 ;
        RECT 146.200 55.100 146.600 55.200 ;
        RECT 147.000 55.100 147.400 59.900 ;
        RECT 149.900 56.300 150.300 59.900 ;
        RECT 149.400 55.900 150.300 56.300 ;
        RECT 146.200 54.800 147.400 55.100 ;
        RECT 145.400 53.800 145.800 54.200 ;
        RECT 145.400 52.100 145.700 53.800 ;
        RECT 145.400 51.100 145.800 52.100 ;
        RECT 147.000 51.100 147.400 54.800 ;
        RECT 149.500 54.200 149.800 55.900 ;
        RECT 150.200 54.800 150.600 55.600 ;
        RECT 149.400 53.800 149.800 54.200 ;
        RECT 147.800 52.400 148.200 53.200 ;
        RECT 148.600 52.400 149.000 53.200 ;
        RECT 149.500 52.200 149.800 53.800 ;
        RECT 149.400 51.100 149.800 52.200 ;
        RECT 0.900 48.400 1.300 49.900 ;
        RECT 0.600 47.900 1.300 48.400 ;
        RECT 3.000 47.900 3.400 49.900 ;
        RECT 5.100 48.200 5.500 49.900 ;
        RECT 6.800 49.200 7.200 49.900 ;
        RECT 10.700 49.200 11.100 49.900 ;
        RECT 6.200 48.800 7.200 49.200 ;
        RECT 10.200 48.800 11.100 49.200 ;
        RECT 4.600 47.900 5.500 48.200 ;
        RECT 0.600 46.200 0.900 47.900 ;
        RECT 3.000 47.800 3.300 47.900 ;
        RECT 2.400 47.600 3.300 47.800 ;
        RECT 1.200 47.500 3.300 47.600 ;
        RECT 1.200 47.300 2.700 47.500 ;
        RECT 1.200 47.200 1.600 47.300 ;
        RECT 0.600 45.800 1.000 46.200 ;
        RECT 0.600 45.100 0.900 45.800 ;
        RECT 1.300 45.500 1.600 47.200 ;
        RECT 2.000 46.600 2.600 47.000 ;
        RECT 2.200 46.200 2.500 46.600 ;
        RECT 3.000 46.400 3.400 47.200 ;
        RECT 3.800 46.800 4.200 47.600 ;
        RECT 2.200 45.800 2.600 46.200 ;
        RECT 4.600 46.100 5.000 47.900 ;
        RECT 5.400 46.800 5.800 47.200 ;
        RECT 6.800 47.100 7.200 48.800 ;
        RECT 10.700 48.200 11.100 48.800 ;
        RECT 10.200 48.100 11.100 48.200 ;
        RECT 11.800 48.100 12.200 48.600 ;
        RECT 10.200 47.800 12.200 48.100 ;
        RECT 6.300 46.900 7.200 47.100 ;
        RECT 6.300 46.800 7.100 46.900 ;
        RECT 9.400 46.800 9.800 47.600 ;
        RECT 5.400 46.100 5.700 46.800 ;
        RECT 4.600 45.800 5.700 46.100 ;
        RECT 1.300 45.200 2.500 45.500 ;
        RECT 0.600 41.100 1.000 45.100 ;
        RECT 2.200 43.100 2.500 45.200 ;
        RECT 2.200 41.100 2.600 43.100 ;
        RECT 4.600 41.100 5.000 45.800 ;
        RECT 6.300 45.200 6.600 46.800 ;
        RECT 7.400 45.800 8.200 46.200 ;
        RECT 5.400 44.400 5.800 45.200 ;
        RECT 6.200 44.800 6.600 45.200 ;
        RECT 8.600 44.800 9.000 45.600 ;
        RECT 6.300 43.500 6.600 44.800 ;
        RECT 7.000 44.100 7.400 44.600 ;
        RECT 7.800 44.100 8.200 44.200 ;
        RECT 7.000 43.800 8.200 44.100 ;
        RECT 6.300 43.200 8.100 43.500 ;
        RECT 6.300 43.100 6.600 43.200 ;
        RECT 6.200 41.100 6.600 43.100 ;
        RECT 7.800 43.100 8.100 43.200 ;
        RECT 7.800 41.100 8.200 43.100 ;
        RECT 10.200 41.100 10.600 47.800 ;
        RECT 12.600 47.100 13.000 49.900 ;
        RECT 13.400 48.000 13.800 49.900 ;
        RECT 15.000 48.000 15.400 49.900 ;
        RECT 13.400 47.900 15.400 48.000 ;
        RECT 15.800 47.900 16.200 49.900 ;
        RECT 17.400 48.900 17.800 49.900 ;
        RECT 13.500 47.700 15.300 47.900 ;
        RECT 13.800 47.200 14.200 47.400 ;
        RECT 15.800 47.200 16.100 47.900 ;
        RECT 16.600 47.800 17.000 48.200 ;
        RECT 13.400 47.100 14.200 47.200 ;
        RECT 12.600 46.900 14.200 47.100 ;
        RECT 12.600 46.800 13.800 46.900 ;
        RECT 14.900 46.800 16.200 47.200 ;
        RECT 16.600 47.100 16.900 47.800 ;
        RECT 17.400 47.200 17.700 48.900 ;
        RECT 18.200 47.800 18.600 48.600 ;
        RECT 19.000 47.900 19.400 49.900 ;
        RECT 21.200 48.100 22.000 49.900 ;
        RECT 19.000 47.600 20.200 47.900 ;
        RECT 19.800 47.500 20.200 47.600 ;
        RECT 20.500 47.400 20.900 47.800 ;
        RECT 20.500 47.200 20.800 47.400 ;
        RECT 17.400 47.100 17.800 47.200 ;
        RECT 16.600 46.800 17.800 47.100 ;
        RECT 19.000 46.800 19.800 47.200 ;
        RECT 20.400 46.800 20.800 47.200 ;
        RECT 11.000 44.400 11.400 45.200 ;
        RECT 12.600 41.100 13.000 46.800 ;
        RECT 14.200 45.800 14.600 46.600 ;
        RECT 14.900 45.200 15.200 46.800 ;
        RECT 16.600 45.400 17.000 46.200 ;
        RECT 14.200 44.800 15.200 45.200 ;
        RECT 15.800 45.100 16.200 45.200 ;
        RECT 17.400 45.100 17.700 46.800 ;
        RECT 21.200 46.400 21.500 48.100 ;
        RECT 23.800 47.900 24.200 49.900 ;
        RECT 24.700 48.200 25.100 48.600 ;
        RECT 21.800 47.700 22.600 47.800 ;
        RECT 21.800 47.400 22.800 47.700 ;
        RECT 23.100 47.600 24.200 47.900 ;
        RECT 24.600 47.800 25.000 48.200 ;
        RECT 25.400 47.900 25.800 49.900 ;
        RECT 27.800 47.900 28.200 49.900 ;
        RECT 28.600 48.000 29.000 49.900 ;
        RECT 30.200 48.000 30.600 49.900 ;
        RECT 28.600 47.900 30.600 48.000 ;
        RECT 31.000 47.900 31.400 49.900 ;
        RECT 31.800 48.000 32.200 49.900 ;
        RECT 33.400 48.000 33.800 49.900 ;
        RECT 31.800 47.900 33.800 48.000 ;
        RECT 34.200 48.000 34.600 49.900 ;
        RECT 35.800 48.000 36.200 49.900 ;
        RECT 34.200 47.900 36.200 48.000 ;
        RECT 36.600 47.900 37.000 49.900 ;
        RECT 37.400 47.900 37.800 49.900 ;
        RECT 38.200 48.000 38.600 49.900 ;
        RECT 39.800 48.000 40.200 49.900 ;
        RECT 38.200 47.900 40.200 48.000 ;
        RECT 41.400 48.900 41.800 49.900 ;
        RECT 23.100 47.500 23.500 47.600 ;
        RECT 22.500 47.200 22.800 47.400 ;
        RECT 21.800 46.700 22.200 47.100 ;
        RECT 22.500 46.900 24.200 47.200 ;
        RECT 23.400 46.800 24.200 46.900 ;
        RECT 21.000 46.200 21.500 46.400 ;
        RECT 20.600 46.100 21.500 46.200 ;
        RECT 21.900 46.400 22.200 46.700 ;
        RECT 21.900 46.100 23.200 46.400 ;
        RECT 20.600 45.800 21.300 46.100 ;
        RECT 22.800 46.000 23.200 46.100 ;
        RECT 24.600 46.100 25.000 46.200 ;
        RECT 25.500 46.100 25.800 47.900 ;
        RECT 27.900 47.200 28.200 47.900 ;
        RECT 28.700 47.700 30.500 47.900 ;
        RECT 29.800 47.200 30.200 47.400 ;
        RECT 31.100 47.200 31.400 47.900 ;
        RECT 31.900 47.700 33.700 47.900 ;
        RECT 34.300 47.700 36.100 47.900 ;
        RECT 33.000 47.200 33.400 47.400 ;
        RECT 34.600 47.200 35.000 47.400 ;
        RECT 36.600 47.200 36.900 47.900 ;
        RECT 37.500 47.200 37.800 47.900 ;
        RECT 38.300 47.700 40.100 47.900 ;
        RECT 39.400 47.200 39.800 47.400 ;
        RECT 41.400 47.200 41.700 48.900 ;
        RECT 42.200 47.800 42.600 48.600 ;
        RECT 43.100 48.200 43.500 48.600 ;
        RECT 43.000 47.800 43.400 48.200 ;
        RECT 43.800 47.900 44.200 49.900 ;
        RECT 46.500 48.200 46.900 49.900 ;
        RECT 50.300 48.200 50.700 48.600 ;
        RECT 26.200 47.100 26.600 47.200 ;
        RECT 27.800 47.100 29.100 47.200 ;
        RECT 26.200 46.800 29.100 47.100 ;
        RECT 29.800 46.900 30.600 47.200 ;
        RECT 30.200 46.800 30.600 46.900 ;
        RECT 31.000 46.800 32.300 47.200 ;
        RECT 33.000 47.100 33.800 47.200 ;
        RECT 34.200 47.100 35.000 47.200 ;
        RECT 33.000 46.900 35.000 47.100 ;
        RECT 33.400 46.800 34.600 46.900 ;
        RECT 35.700 46.800 37.000 47.200 ;
        RECT 37.400 46.800 38.700 47.200 ;
        RECT 39.400 46.900 40.200 47.200 ;
        RECT 39.800 46.800 40.200 46.900 ;
        RECT 41.400 46.800 41.800 47.200 ;
        RECT 43.000 47.100 43.400 47.200 ;
        RECT 43.900 47.100 44.200 47.900 ;
        RECT 43.000 46.800 44.200 47.100 ;
        RECT 46.200 47.800 47.400 48.200 ;
        RECT 50.200 47.800 50.600 48.200 ;
        RECT 51.000 47.900 51.400 49.900 ;
        RECT 53.700 49.200 54.100 49.900 ;
        RECT 53.400 48.800 54.100 49.200 ;
        RECT 53.700 48.200 54.100 48.800 ;
        RECT 57.100 49.200 57.500 49.900 ;
        RECT 57.100 48.800 57.800 49.200 ;
        RECT 57.100 48.200 57.500 48.800 ;
        RECT 53.700 47.900 54.600 48.200 ;
        RECT 46.200 47.200 46.500 47.800 ;
        RECT 46.200 46.800 46.600 47.200 ;
        RECT 26.200 46.400 26.600 46.800 ;
        RECT 27.000 46.100 27.400 46.200 ;
        RECT 24.600 45.800 25.800 46.100 ;
        RECT 26.600 45.800 27.400 46.100 ;
        RECT 21.000 45.100 21.300 45.800 ;
        RECT 21.700 45.700 22.100 45.800 ;
        RECT 21.700 45.400 23.400 45.700 ;
        RECT 23.100 45.100 23.400 45.400 ;
        RECT 24.700 45.100 25.000 45.800 ;
        RECT 26.600 45.600 27.000 45.800 ;
        RECT 27.800 45.100 28.200 45.200 ;
        RECT 28.800 45.100 29.100 46.800 ;
        RECT 29.400 45.800 29.800 46.600 ;
        RECT 31.000 45.100 31.400 45.200 ;
        RECT 32.000 45.100 32.300 46.800 ;
        RECT 32.600 46.100 33.000 46.600 ;
        RECT 35.000 46.100 35.400 46.600 ;
        RECT 32.600 45.800 35.400 46.100 ;
        RECT 35.700 45.100 36.000 46.800 ;
        RECT 36.600 45.100 37.000 45.200 ;
        RECT 37.400 45.100 37.800 45.200 ;
        RECT 38.400 45.100 38.700 46.800 ;
        RECT 39.000 45.800 39.400 46.600 ;
        RECT 40.600 45.400 41.000 46.200 ;
        RECT 41.400 45.100 41.700 46.800 ;
        RECT 43.000 46.100 43.400 46.200 ;
        RECT 43.900 46.100 44.200 46.800 ;
        RECT 45.400 46.100 45.800 46.200 ;
        RECT 43.000 45.800 44.200 46.100 ;
        RECT 45.000 45.800 45.800 46.100 ;
        RECT 43.100 45.100 43.400 45.800 ;
        RECT 45.000 45.600 45.400 45.800 ;
        RECT 15.500 44.800 16.200 45.100 ;
        RECT 14.700 41.100 15.100 44.800 ;
        RECT 15.500 44.200 15.800 44.800 ;
        RECT 15.400 43.800 15.800 44.200 ;
        RECT 16.900 44.700 17.800 45.100 ;
        RECT 19.000 44.800 20.200 45.100 ;
        RECT 21.000 44.800 22.000 45.100 ;
        RECT 16.900 41.100 17.300 44.700 ;
        RECT 19.000 41.100 19.400 44.800 ;
        RECT 19.800 44.700 20.200 44.800 ;
        RECT 21.200 41.100 22.000 44.800 ;
        RECT 23.100 44.800 24.200 45.100 ;
        RECT 23.100 44.700 23.500 44.800 ;
        RECT 23.800 41.100 24.200 44.800 ;
        RECT 24.600 41.100 25.000 45.100 ;
        RECT 25.400 44.800 27.400 45.100 ;
        RECT 27.800 44.800 28.500 45.100 ;
        RECT 28.800 44.800 29.300 45.100 ;
        RECT 31.000 44.800 31.700 45.100 ;
        RECT 32.000 44.800 32.500 45.100 ;
        RECT 25.400 41.100 25.800 44.800 ;
        RECT 27.000 41.100 27.400 44.800 ;
        RECT 28.200 44.200 28.500 44.800 ;
        RECT 28.200 43.800 28.600 44.200 ;
        RECT 28.900 41.100 29.300 44.800 ;
        RECT 31.400 44.200 31.700 44.800 ;
        RECT 31.400 43.800 31.800 44.200 ;
        RECT 32.100 41.100 32.500 44.800 ;
        RECT 35.500 44.800 36.000 45.100 ;
        RECT 36.300 44.800 38.100 45.100 ;
        RECT 38.400 44.800 38.900 45.100 ;
        RECT 35.500 41.100 35.900 44.800 ;
        RECT 36.300 44.200 36.600 44.800 ;
        RECT 36.200 43.800 36.600 44.200 ;
        RECT 37.800 44.200 38.100 44.800 ;
        RECT 37.800 43.800 38.200 44.200 ;
        RECT 38.500 41.100 38.900 44.800 ;
        RECT 40.900 44.700 41.800 45.100 ;
        RECT 40.900 44.200 41.300 44.700 ;
        RECT 40.600 43.800 41.300 44.200 ;
        RECT 40.900 41.100 41.300 43.800 ;
        RECT 43.000 41.100 43.400 45.100 ;
        RECT 43.800 44.800 45.800 45.100 ;
        RECT 43.800 41.100 44.200 44.800 ;
        RECT 45.400 41.100 45.800 44.800 ;
        RECT 47.000 41.100 47.400 47.800 ;
        RECT 47.800 46.800 48.200 47.600 ;
        RECT 49.400 47.100 49.800 47.200 ;
        RECT 51.100 47.100 51.400 47.900 ;
        RECT 49.400 46.800 51.400 47.100 ;
        RECT 50.200 46.100 50.600 46.200 ;
        RECT 51.100 46.100 51.400 46.800 ;
        RECT 52.600 46.100 53.000 46.200 ;
        RECT 50.200 45.800 51.400 46.100 ;
        RECT 52.200 45.800 53.000 46.100 ;
        RECT 50.300 45.100 50.600 45.800 ;
        RECT 52.200 45.600 52.600 45.800 ;
        RECT 50.200 41.100 50.600 45.100 ;
        RECT 51.000 44.800 53.000 45.100 ;
        RECT 51.000 41.100 51.400 44.800 ;
        RECT 52.600 41.100 53.000 44.800 ;
        RECT 54.200 41.100 54.600 47.900 ;
        RECT 56.600 47.900 57.500 48.200 ;
        RECT 58.200 47.900 58.600 49.900 ;
        RECT 59.000 48.000 59.400 49.900 ;
        RECT 60.600 48.000 61.000 49.900 ;
        RECT 61.700 49.200 62.100 49.900 ;
        RECT 61.400 48.800 62.100 49.200 ;
        RECT 59.000 47.900 61.000 48.000 ;
        RECT 61.700 48.200 62.100 48.800 ;
        RECT 64.600 48.200 65.000 49.900 ;
        RECT 61.700 47.900 62.600 48.200 ;
        RECT 55.000 46.800 55.400 47.600 ;
        RECT 55.800 46.800 56.200 47.600 ;
        RECT 56.600 41.100 57.000 47.900 ;
        RECT 58.300 47.200 58.600 47.900 ;
        RECT 59.100 47.700 60.900 47.900 ;
        RECT 60.200 47.200 60.600 47.400 ;
        RECT 57.400 47.100 57.800 47.200 ;
        RECT 58.200 47.100 59.500 47.200 ;
        RECT 57.400 46.800 59.500 47.100 ;
        RECT 60.200 46.900 61.000 47.200 ;
        RECT 60.600 46.800 61.000 46.900 ;
        RECT 58.200 45.100 58.600 45.200 ;
        RECT 59.200 45.100 59.500 46.800 ;
        RECT 59.800 45.800 60.200 46.600 ;
        RECT 58.200 44.800 58.900 45.100 ;
        RECT 59.200 44.800 59.700 45.100 ;
        RECT 58.600 44.200 58.900 44.800 ;
        RECT 58.600 43.800 59.000 44.200 ;
        RECT 59.300 41.100 59.700 44.800 ;
        RECT 62.200 41.100 62.600 47.900 ;
        RECT 64.500 47.900 65.000 48.200 ;
        RECT 63.000 47.100 63.400 47.600 ;
        RECT 64.500 47.200 64.800 47.900 ;
        RECT 66.200 47.600 66.600 49.900 ;
        RECT 65.300 47.300 66.600 47.600 ;
        RECT 67.000 47.600 67.400 49.900 ;
        RECT 68.600 48.200 69.000 49.900 ;
        RECT 70.500 49.200 70.900 49.900 ;
        RECT 70.200 48.800 70.900 49.200 ;
        RECT 70.500 48.200 70.900 48.800 ;
        RECT 72.900 48.200 73.300 49.900 ;
        RECT 68.600 47.900 69.100 48.200 ;
        RECT 70.500 47.900 71.400 48.200 ;
        RECT 67.000 47.300 68.300 47.600 ;
        RECT 64.500 47.100 65.000 47.200 ;
        RECT 63.000 46.800 65.000 47.100 ;
        RECT 64.500 45.100 64.800 46.800 ;
        RECT 65.300 46.500 65.600 47.300 ;
        RECT 65.100 46.100 65.600 46.500 ;
        RECT 65.300 45.100 65.600 46.100 ;
        RECT 68.000 46.500 68.300 47.300 ;
        RECT 68.800 47.200 69.100 47.900 ;
        RECT 68.600 47.100 69.100 47.200 ;
        RECT 70.200 47.100 70.600 47.200 ;
        RECT 68.600 46.800 70.600 47.100 ;
        RECT 68.000 46.100 68.500 46.500 ;
        RECT 68.000 45.100 68.300 46.100 ;
        RECT 68.800 45.100 69.100 46.800 ;
        RECT 64.500 44.600 65.000 45.100 ;
        RECT 65.300 44.800 66.600 45.100 ;
        RECT 64.600 41.100 65.000 44.600 ;
        RECT 66.200 41.100 66.600 44.800 ;
        RECT 67.000 44.800 68.300 45.100 ;
        RECT 67.000 41.100 67.400 44.800 ;
        RECT 68.600 44.600 69.100 45.100 ;
        RECT 68.600 41.100 69.000 44.600 ;
        RECT 71.000 41.100 71.400 47.900 ;
        RECT 72.600 47.800 73.800 48.200 ;
        RECT 75.000 47.900 75.400 49.900 ;
        RECT 75.800 48.000 76.200 49.900 ;
        RECT 77.400 48.000 77.800 49.900 ;
        RECT 75.800 47.900 77.800 48.000 ;
        RECT 79.000 48.900 79.400 49.900 ;
        RECT 71.800 46.800 72.200 47.600 ;
        RECT 72.600 47.200 72.900 47.800 ;
        RECT 72.600 46.800 73.000 47.200 ;
        RECT 73.400 41.100 73.800 47.800 ;
        RECT 74.200 46.800 74.600 47.600 ;
        RECT 75.100 47.200 75.400 47.900 ;
        RECT 75.900 47.700 77.700 47.900 ;
        RECT 77.000 47.200 77.400 47.400 ;
        RECT 79.000 47.200 79.300 48.900 ;
        RECT 79.800 47.800 80.200 48.600 ;
        RECT 80.600 48.000 81.000 49.900 ;
        RECT 82.200 48.000 82.600 49.900 ;
        RECT 80.600 47.900 82.600 48.000 ;
        RECT 83.000 47.900 83.400 49.900 ;
        RECT 83.800 48.000 84.200 49.900 ;
        RECT 85.400 48.000 85.800 49.900 ;
        RECT 83.800 47.900 85.800 48.000 ;
        RECT 86.200 47.900 86.600 49.900 ;
        RECT 87.000 47.900 87.400 49.900 ;
        RECT 87.800 48.000 88.200 49.900 ;
        RECT 89.400 48.000 89.800 49.900 ;
        RECT 87.800 47.900 89.800 48.000 ;
        RECT 90.200 48.000 90.600 49.900 ;
        RECT 91.800 48.000 92.200 49.900 ;
        RECT 90.200 47.900 92.200 48.000 ;
        RECT 92.600 47.900 93.000 49.900 ;
        RECT 93.700 48.200 94.100 49.900 ;
        RECT 93.700 47.900 94.600 48.200 ;
        RECT 95.800 48.000 96.200 49.900 ;
        RECT 97.400 48.000 97.800 49.900 ;
        RECT 95.800 47.900 97.800 48.000 ;
        RECT 98.200 47.900 98.600 49.900 ;
        RECT 100.600 49.600 102.600 49.900 ;
        RECT 100.600 47.900 101.000 49.600 ;
        RECT 101.400 47.900 101.800 49.300 ;
        RECT 102.200 48.000 102.600 49.600 ;
        RECT 103.800 48.000 104.200 49.900 ;
        RECT 102.200 47.900 104.200 48.000 ;
        RECT 104.600 47.900 105.000 49.900 ;
        RECT 105.400 48.000 105.800 49.900 ;
        RECT 107.000 48.000 107.400 49.900 ;
        RECT 105.400 47.900 107.400 48.000 ;
        RECT 107.800 48.000 108.200 49.900 ;
        RECT 109.400 48.000 109.800 49.900 ;
        RECT 107.800 47.900 109.800 48.000 ;
        RECT 110.200 47.900 110.600 49.900 ;
        RECT 80.700 47.700 82.500 47.900 ;
        RECT 81.000 47.200 81.400 47.400 ;
        RECT 83.000 47.200 83.300 47.900 ;
        RECT 83.900 47.700 85.700 47.900 ;
        RECT 84.200 47.200 84.600 47.400 ;
        RECT 86.200 47.200 86.500 47.900 ;
        RECT 87.100 47.200 87.400 47.900 ;
        RECT 87.900 47.700 89.700 47.900 ;
        RECT 90.300 47.700 92.100 47.900 ;
        RECT 89.000 47.200 89.400 47.400 ;
        RECT 90.600 47.200 91.000 47.400 ;
        RECT 92.600 47.200 92.900 47.900 ;
        RECT 75.000 46.800 76.300 47.200 ;
        RECT 77.000 46.900 77.800 47.200 ;
        RECT 77.400 46.800 77.800 46.900 ;
        RECT 79.000 46.800 79.400 47.200 ;
        RECT 80.600 46.900 81.400 47.200 ;
        RECT 80.600 46.800 81.000 46.900 ;
        RECT 82.100 46.800 83.400 47.200 ;
        RECT 83.800 46.900 84.600 47.200 ;
        RECT 83.800 46.800 84.200 46.900 ;
        RECT 85.300 46.800 86.600 47.200 ;
        RECT 87.000 46.800 88.300 47.200 ;
        RECT 89.000 46.900 89.800 47.200 ;
        RECT 89.400 46.800 89.800 46.900 ;
        RECT 90.200 46.900 91.000 47.200 ;
        RECT 91.700 47.100 93.000 47.200 ;
        RECT 93.400 47.100 93.800 47.200 ;
        RECT 90.200 46.800 90.600 46.900 ;
        RECT 91.700 46.800 93.800 47.100 ;
        RECT 74.200 45.100 74.600 45.200 ;
        RECT 75.000 45.100 75.400 45.200 ;
        RECT 76.000 45.100 76.300 46.800 ;
        RECT 76.600 45.800 77.000 46.600 ;
        RECT 79.000 46.200 79.300 46.800 ;
        RECT 78.200 45.400 78.600 46.200 ;
        RECT 79.000 45.800 79.400 46.200 ;
        RECT 81.400 45.800 81.800 46.600 ;
        RECT 79.000 45.100 79.300 45.800 ;
        RECT 82.100 45.100 82.400 46.800 ;
        RECT 83.000 46.100 83.400 46.200 ;
        RECT 84.600 46.100 85.000 46.600 ;
        RECT 83.000 45.800 85.000 46.100 ;
        RECT 85.300 46.200 85.600 46.800 ;
        RECT 85.300 45.800 85.800 46.200 ;
        RECT 83.000 45.100 83.400 45.200 ;
        RECT 85.300 45.100 85.600 45.800 ;
        RECT 86.200 45.100 86.600 45.200 ;
        RECT 74.200 44.800 75.700 45.100 ;
        RECT 76.000 44.800 76.500 45.100 ;
        RECT 75.400 44.200 75.700 44.800 ;
        RECT 75.400 43.800 75.800 44.200 ;
        RECT 76.100 42.200 76.500 44.800 ;
        RECT 78.500 44.700 79.400 45.100 ;
        RECT 81.900 44.800 82.400 45.100 ;
        RECT 82.700 44.800 83.400 45.100 ;
        RECT 85.100 44.800 85.600 45.100 ;
        RECT 85.900 44.800 86.600 45.100 ;
        RECT 87.000 45.100 87.400 45.200 ;
        RECT 88.000 45.100 88.300 46.800 ;
        RECT 88.600 45.800 89.000 46.600 ;
        RECT 91.000 45.800 91.400 46.600 ;
        RECT 91.700 45.100 92.000 46.800 ;
        RECT 94.200 46.100 94.600 47.900 ;
        RECT 95.900 47.700 97.700 47.900 ;
        RECT 92.600 45.800 94.600 46.100 ;
        RECT 92.600 45.200 92.900 45.800 ;
        RECT 92.600 45.100 93.000 45.200 ;
        RECT 87.000 44.800 87.700 45.100 ;
        RECT 88.000 44.800 88.500 45.100 ;
        RECT 76.100 41.800 77.000 42.200 ;
        RECT 76.100 41.100 76.500 41.800 ;
        RECT 78.500 41.100 78.900 44.700 ;
        RECT 81.900 41.100 82.300 44.800 ;
        RECT 82.700 44.200 83.000 44.800 ;
        RECT 82.600 43.800 83.000 44.200 ;
        RECT 85.100 41.100 85.500 44.800 ;
        RECT 85.900 44.200 86.200 44.800 ;
        RECT 85.800 43.800 86.200 44.200 ;
        RECT 87.400 44.200 87.700 44.800 ;
        RECT 87.400 43.800 87.800 44.200 ;
        RECT 88.100 41.100 88.500 44.800 ;
        RECT 91.500 44.800 92.000 45.100 ;
        RECT 92.300 44.800 93.000 45.100 ;
        RECT 91.500 41.100 91.900 44.800 ;
        RECT 92.300 44.200 92.600 44.800 ;
        RECT 93.400 44.400 93.800 45.200 ;
        RECT 92.200 43.800 92.600 44.200 ;
        RECT 94.200 41.100 94.600 45.800 ;
        RECT 95.000 46.800 95.400 47.600 ;
        RECT 96.200 47.200 96.600 47.400 ;
        RECT 98.200 47.200 98.500 47.900 ;
        RECT 101.400 47.200 101.700 47.900 ;
        RECT 102.300 47.700 104.100 47.900 ;
        RECT 103.400 47.200 103.800 47.400 ;
        RECT 104.700 47.200 105.000 47.900 ;
        RECT 105.500 47.700 107.300 47.900 ;
        RECT 107.900 47.700 109.700 47.900 ;
        RECT 106.600 47.200 107.000 47.400 ;
        RECT 108.200 47.200 108.600 47.400 ;
        RECT 110.200 47.200 110.500 47.900 ;
        RECT 95.800 46.900 96.600 47.200 ;
        RECT 95.800 46.800 96.200 46.900 ;
        RECT 97.300 46.800 98.600 47.200 ;
        RECT 95.000 46.100 95.300 46.800 ;
        RECT 96.600 46.100 97.000 46.600 ;
        RECT 95.000 45.800 97.000 46.100 ;
        RECT 97.300 46.100 97.600 46.800 ;
        RECT 100.600 46.400 101.000 47.200 ;
        RECT 101.400 46.900 102.600 47.200 ;
        RECT 103.400 46.900 104.200 47.200 ;
        RECT 102.200 46.800 102.600 46.900 ;
        RECT 103.800 46.800 104.200 46.900 ;
        RECT 104.600 46.800 105.900 47.200 ;
        RECT 106.600 46.900 107.400 47.200 ;
        RECT 107.000 46.800 107.400 46.900 ;
        RECT 107.800 46.900 108.600 47.200 ;
        RECT 107.800 46.800 108.200 46.900 ;
        RECT 109.300 46.800 110.600 47.200 ;
        RECT 99.800 46.100 100.200 46.200 ;
        RECT 97.300 45.800 100.200 46.100 ;
        RECT 101.400 45.800 101.800 46.600 ;
        RECT 95.000 45.200 95.300 45.800 ;
        RECT 95.000 44.800 95.400 45.200 ;
        RECT 97.300 45.100 97.600 45.800 ;
        RECT 98.200 45.100 98.600 45.200 ;
        RECT 99.000 45.100 99.400 45.200 ;
        RECT 102.300 45.100 102.600 46.800 ;
        RECT 103.000 45.800 103.400 46.600 ;
        RECT 104.600 45.100 105.000 45.200 ;
        RECT 105.600 45.100 105.900 46.800 ;
        RECT 106.200 45.800 106.600 46.600 ;
        RECT 108.600 45.800 109.000 46.600 ;
        RECT 109.300 45.100 109.600 46.800 ;
        RECT 110.200 45.100 110.600 45.200 ;
        RECT 97.100 44.800 97.600 45.100 ;
        RECT 97.900 44.800 99.400 45.100 ;
        RECT 97.100 41.100 97.500 44.800 ;
        RECT 97.900 44.200 98.200 44.800 ;
        RECT 97.800 43.800 98.200 44.200 ;
        RECT 101.900 41.100 102.900 45.100 ;
        RECT 104.600 44.800 105.300 45.100 ;
        RECT 105.600 44.800 106.100 45.100 ;
        RECT 105.000 44.200 105.300 44.800 ;
        RECT 105.000 43.800 105.400 44.200 ;
        RECT 105.700 41.100 106.100 44.800 ;
        RECT 109.100 44.800 109.600 45.100 ;
        RECT 109.900 44.800 110.600 45.100 ;
        RECT 109.100 42.200 109.500 44.800 ;
        RECT 109.900 44.200 110.200 44.800 ;
        RECT 109.800 43.800 110.200 44.200 ;
        RECT 108.600 41.800 109.500 42.200 ;
        RECT 109.100 41.100 109.500 41.800 ;
        RECT 111.000 41.100 111.400 49.900 ;
        RECT 113.400 48.800 113.800 49.900 ;
        RECT 111.800 47.800 112.200 48.600 ;
        RECT 112.600 47.800 113.000 48.600 ;
        RECT 113.500 47.200 113.800 48.800 ;
        RECT 115.000 48.000 115.400 49.900 ;
        RECT 116.600 48.000 117.000 49.900 ;
        RECT 115.000 47.900 117.000 48.000 ;
        RECT 117.400 47.900 117.800 49.900 ;
        RECT 118.200 48.000 118.600 49.900 ;
        RECT 119.800 48.000 120.200 49.900 ;
        RECT 118.200 47.900 120.200 48.000 ;
        RECT 120.600 47.900 121.000 49.900 ;
        RECT 121.700 48.200 122.100 49.900 ;
        RECT 121.700 47.900 122.600 48.200 ;
        RECT 115.100 47.700 116.900 47.900 ;
        RECT 115.400 47.200 115.800 47.400 ;
        RECT 117.400 47.200 117.700 47.900 ;
        RECT 118.300 47.700 120.100 47.900 ;
        RECT 118.600 47.200 119.000 47.400 ;
        RECT 120.600 47.200 120.900 47.900 ;
        RECT 113.400 47.100 113.800 47.200 ;
        RECT 115.000 47.100 115.800 47.200 ;
        RECT 113.400 46.900 115.800 47.100 ;
        RECT 113.400 46.800 115.400 46.900 ;
        RECT 116.500 46.800 117.800 47.200 ;
        RECT 118.200 46.900 119.000 47.200 ;
        RECT 118.200 46.800 118.600 46.900 ;
        RECT 119.700 46.800 121.000 47.200 ;
        RECT 113.500 45.100 113.800 46.800 ;
        RECT 114.200 46.100 114.600 46.200 ;
        RECT 115.000 46.100 115.400 46.200 ;
        RECT 114.200 45.800 115.400 46.100 ;
        RECT 115.800 45.800 116.200 46.600 ;
        RECT 114.200 45.400 114.600 45.800 ;
        RECT 116.500 45.100 116.800 46.800 ;
        RECT 119.000 45.800 119.400 46.600 ;
        RECT 117.400 45.100 117.800 45.200 ;
        RECT 119.700 45.100 120.000 46.800 ;
        RECT 121.400 46.100 121.800 46.200 ;
        RECT 122.200 46.100 122.600 47.900 ;
        RECT 125.400 47.900 125.800 49.900 ;
        RECT 126.100 48.200 126.500 48.600 ;
        RECT 123.000 46.800 123.400 47.600 ;
        RECT 124.600 46.400 125.000 47.200 ;
        RECT 121.400 45.800 122.600 46.100 ;
        RECT 123.800 46.100 124.200 46.200 ;
        RECT 125.400 46.100 125.700 47.900 ;
        RECT 126.200 47.800 126.600 48.200 ;
        RECT 127.000 47.900 127.400 49.900 ;
        RECT 127.800 48.000 128.200 49.900 ;
        RECT 129.400 48.000 129.800 49.900 ;
        RECT 127.800 47.900 129.800 48.000 ;
        RECT 127.100 47.200 127.400 47.900 ;
        RECT 127.900 47.700 129.700 47.900 ;
        RECT 129.000 47.200 129.400 47.400 ;
        RECT 126.200 47.100 126.600 47.200 ;
        RECT 127.000 47.100 128.300 47.200 ;
        RECT 126.200 46.800 128.300 47.100 ;
        RECT 129.000 46.900 129.800 47.200 ;
        RECT 132.000 47.100 132.400 49.900 ;
        RECT 132.000 46.900 132.900 47.100 ;
        RECT 129.400 46.800 129.800 46.900 ;
        RECT 132.100 46.800 132.900 46.900 ;
        RECT 126.200 46.100 126.600 46.200 ;
        RECT 127.000 46.100 127.400 46.200 ;
        RECT 123.800 45.800 124.600 46.100 ;
        RECT 125.400 45.800 127.400 46.100 ;
        RECT 120.600 45.100 121.000 45.200 ;
        RECT 113.400 44.700 114.300 45.100 ;
        RECT 113.900 41.100 114.300 44.700 ;
        RECT 116.300 44.800 116.800 45.100 ;
        RECT 117.100 44.800 117.800 45.100 ;
        RECT 119.500 44.800 120.000 45.100 ;
        RECT 120.300 44.800 121.000 45.100 ;
        RECT 116.300 42.200 116.700 44.800 ;
        RECT 117.100 44.200 117.400 44.800 ;
        RECT 117.000 43.800 117.400 44.200 ;
        RECT 115.800 41.800 116.700 42.200 ;
        RECT 116.300 41.100 116.700 41.800 ;
        RECT 119.500 41.100 119.900 44.800 ;
        RECT 120.300 44.200 120.600 44.800 ;
        RECT 121.400 44.400 121.800 45.200 ;
        RECT 120.200 43.800 120.600 44.200 ;
        RECT 122.200 41.100 122.600 45.800 ;
        RECT 124.200 45.600 124.600 45.800 ;
        RECT 126.200 45.100 126.500 45.800 ;
        RECT 128.000 45.100 128.300 46.800 ;
        RECT 128.600 45.800 129.000 46.600 ;
        RECT 131.000 45.800 131.800 46.200 ;
        RECT 123.800 44.800 125.800 45.100 ;
        RECT 123.800 41.100 124.200 44.800 ;
        RECT 125.400 41.100 125.800 44.800 ;
        RECT 126.200 41.100 126.600 45.100 ;
        RECT 128.000 44.800 128.500 45.100 ;
        RECT 130.200 44.800 130.600 45.600 ;
        RECT 132.600 45.200 132.900 46.800 ;
        RECT 128.100 41.100 128.500 44.800 ;
        RECT 131.800 43.800 132.200 45.200 ;
        RECT 132.600 44.800 133.000 45.200 ;
        RECT 132.600 43.500 132.900 44.800 ;
        RECT 131.100 43.200 132.900 43.500 ;
        RECT 131.100 43.100 131.400 43.200 ;
        RECT 131.000 41.100 131.400 43.100 ;
        RECT 132.600 43.100 132.900 43.200 ;
        RECT 132.600 41.100 133.000 43.100 ;
        RECT 133.400 41.100 133.800 49.900 ;
        RECT 135.800 48.900 136.200 49.900 ;
        RECT 135.000 47.800 135.400 48.600 ;
        RECT 134.200 46.800 134.600 47.600 ;
        RECT 135.900 47.200 136.200 48.900 ;
        RECT 135.800 46.800 136.200 47.200 ;
        RECT 135.900 45.100 136.200 46.800 ;
        RECT 136.600 45.400 137.000 46.200 ;
        RECT 135.800 44.700 136.700 45.100 ;
        RECT 136.300 44.200 136.700 44.700 ;
        RECT 136.300 43.800 137.000 44.200 ;
        RECT 136.300 41.100 136.700 43.800 ;
        RECT 138.200 41.100 138.600 49.900 ;
        RECT 141.400 47.900 141.800 49.900 ;
        RECT 142.100 48.200 142.500 48.600 ;
        RECT 143.300 48.200 143.700 49.900 ;
        RECT 142.200 48.100 142.600 48.200 ;
        RECT 143.300 48.100 144.200 48.200 ;
        RECT 139.000 47.100 139.400 47.600 ;
        RECT 139.800 47.100 140.200 47.200 ;
        RECT 139.000 46.800 140.200 47.100 ;
        RECT 140.600 46.400 141.000 47.200 ;
        RECT 139.800 46.100 140.200 46.200 ;
        RECT 141.400 46.100 141.700 47.900 ;
        RECT 142.200 47.800 144.200 48.100 ;
        RECT 145.400 47.900 145.800 49.900 ;
        RECT 146.200 48.000 146.600 49.900 ;
        RECT 147.800 48.000 148.200 49.900 ;
        RECT 149.400 48.800 149.800 49.900 ;
        RECT 146.200 47.900 148.200 48.000 ;
        RECT 142.200 46.100 142.600 46.200 ;
        RECT 139.800 45.800 140.600 46.100 ;
        RECT 141.400 45.800 142.600 46.100 ;
        RECT 140.200 45.600 140.600 45.800 ;
        RECT 142.200 45.100 142.500 45.800 ;
        RECT 139.800 44.800 141.800 45.100 ;
        RECT 139.800 41.100 140.200 44.800 ;
        RECT 141.400 41.100 141.800 44.800 ;
        RECT 142.200 41.100 142.600 45.100 ;
        RECT 143.000 44.400 143.400 45.200 ;
        RECT 143.800 41.100 144.200 47.800 ;
        RECT 144.600 47.100 145.000 47.600 ;
        RECT 145.500 47.200 145.800 47.900 ;
        RECT 146.300 47.700 148.100 47.900 ;
        RECT 147.400 47.200 147.800 47.400 ;
        RECT 149.500 47.200 149.800 48.800 ;
        RECT 145.400 47.100 146.700 47.200 ;
        RECT 144.600 46.800 146.700 47.100 ;
        RECT 147.400 46.900 148.200 47.200 ;
        RECT 147.800 46.800 148.200 46.900 ;
        RECT 149.400 46.800 149.800 47.200 ;
        RECT 145.400 45.100 145.800 45.200 ;
        RECT 146.400 45.100 146.700 46.800 ;
        RECT 147.000 46.100 147.400 46.600 ;
        RECT 149.500 46.100 149.800 46.800 ;
        RECT 147.000 45.800 149.800 46.100 ;
        RECT 149.500 45.100 149.800 45.800 ;
        RECT 150.200 45.400 150.600 46.200 ;
        RECT 145.400 44.800 146.100 45.100 ;
        RECT 146.400 44.800 146.900 45.100 ;
        RECT 145.800 44.200 146.100 44.800 ;
        RECT 145.800 43.800 146.200 44.200 ;
        RECT 146.500 41.100 146.900 44.800 ;
        RECT 149.400 44.700 150.300 45.100 ;
        RECT 149.900 41.100 150.300 44.700 ;
        RECT 1.700 39.200 2.100 39.900 ;
        RECT 1.700 38.800 2.600 39.200 ;
        RECT 1.000 36.800 1.400 37.200 ;
        RECT 1.000 36.200 1.300 36.800 ;
        RECT 1.700 36.200 2.100 38.800 ;
        RECT 0.600 35.900 1.300 36.200 ;
        RECT 1.600 35.900 2.100 36.200 ;
        RECT 3.800 36.200 4.200 39.900 ;
        RECT 5.400 36.200 5.800 39.900 ;
        RECT 3.800 35.900 5.800 36.200 ;
        RECT 6.200 35.900 6.600 39.900 ;
        RECT 7.800 37.900 8.200 39.900 ;
        RECT 7.900 37.800 8.200 37.900 ;
        RECT 9.400 37.900 9.800 39.900 ;
        RECT 11.500 39.200 11.900 39.900 ;
        RECT 11.000 38.800 11.900 39.200 ;
        RECT 9.400 37.800 9.700 37.900 ;
        RECT 7.900 37.500 9.700 37.800 ;
        RECT 8.600 36.400 9.000 37.200 ;
        RECT 9.400 36.200 9.700 37.500 ;
        RECT 11.500 36.200 11.900 38.800 ;
        RECT 14.200 37.900 14.600 39.900 ;
        RECT 14.300 37.800 14.600 37.900 ;
        RECT 15.800 37.900 16.200 39.900 ;
        RECT 15.800 37.800 16.100 37.900 ;
        RECT 14.300 37.500 16.100 37.800 ;
        RECT 12.200 36.800 12.600 37.200 ;
        RECT 12.300 36.200 12.600 36.800 ;
        RECT 15.000 36.400 15.400 37.200 ;
        RECT 15.800 36.200 16.100 37.500 ;
        RECT 0.600 35.800 1.000 35.900 ;
        RECT 1.600 34.200 1.900 35.900 ;
        RECT 4.200 35.200 4.600 35.400 ;
        RECT 6.200 35.200 6.500 35.900 ;
        RECT 7.000 35.400 7.400 36.200 ;
        RECT 9.400 35.800 9.800 36.200 ;
        RECT 11.500 35.900 12.000 36.200 ;
        RECT 12.300 35.900 13.000 36.200 ;
        RECT 2.200 34.400 2.600 35.200 ;
        RECT 3.800 34.900 4.600 35.200 ;
        RECT 5.400 34.900 6.600 35.200 ;
        RECT 3.800 34.800 4.200 34.900 ;
        RECT 0.600 33.800 1.900 34.200 ;
        RECT 3.000 34.100 3.400 34.200 ;
        RECT 2.600 33.800 3.400 34.100 ;
        RECT 4.600 33.800 5.000 34.600 ;
        RECT 5.400 34.200 5.700 34.900 ;
        RECT 6.200 34.800 6.600 34.900 ;
        RECT 7.800 34.800 8.600 35.200 ;
        RECT 9.400 34.200 9.700 35.800 ;
        RECT 11.000 34.400 11.400 35.200 ;
        RECT 11.700 34.200 12.000 35.900 ;
        RECT 12.600 35.800 13.000 35.900 ;
        RECT 13.400 35.400 13.800 36.200 ;
        RECT 15.800 35.800 16.200 36.200 ;
        RECT 16.600 35.900 17.000 39.900 ;
        RECT 17.400 36.200 17.800 39.900 ;
        RECT 19.000 36.200 19.400 39.900 ;
        RECT 20.600 37.900 21.000 39.900 ;
        RECT 20.700 37.800 21.000 37.900 ;
        RECT 22.200 37.900 22.600 39.900 ;
        RECT 22.200 37.800 22.500 37.900 ;
        RECT 20.700 37.500 22.500 37.800 ;
        RECT 21.400 36.400 21.800 37.200 ;
        RECT 22.200 36.200 22.500 37.500 ;
        RECT 23.000 36.200 23.400 39.900 ;
        RECT 23.900 36.200 24.300 36.300 ;
        RECT 25.200 36.200 26.000 39.900 ;
        RECT 17.400 35.900 19.400 36.200 ;
        RECT 14.200 34.800 15.000 35.200 ;
        RECT 15.800 34.200 16.100 35.800 ;
        RECT 16.700 35.200 17.000 35.900 ;
        RECT 18.600 35.200 19.000 35.400 ;
        RECT 5.400 33.800 5.800 34.200 ;
        RECT 8.900 34.100 9.700 34.200 ;
        RECT 8.800 33.900 9.700 34.100 ;
        RECT 10.200 34.100 10.600 34.200 ;
        RECT 0.700 33.100 1.000 33.800 ;
        RECT 2.600 33.600 3.000 33.800 ;
        RECT 1.500 33.100 3.300 33.300 ;
        RECT 5.400 33.100 5.700 33.800 ;
        RECT 0.600 31.100 1.000 33.100 ;
        RECT 1.400 33.000 3.400 33.100 ;
        RECT 1.400 31.100 1.800 33.000 ;
        RECT 3.000 31.100 3.400 33.000 ;
        RECT 5.400 31.100 5.800 33.100 ;
        RECT 6.200 32.800 6.600 33.200 ;
        RECT 6.100 32.400 6.500 32.800 ;
        RECT 8.800 31.100 9.200 33.900 ;
        RECT 10.200 33.800 11.000 34.100 ;
        RECT 11.700 33.800 13.000 34.200 ;
        RECT 15.300 34.100 16.100 34.200 ;
        RECT 15.200 33.900 16.100 34.100 ;
        RECT 16.600 34.900 17.800 35.200 ;
        RECT 18.600 35.100 19.400 35.200 ;
        RECT 19.800 35.100 20.200 36.200 ;
        RECT 22.200 35.800 22.600 36.200 ;
        RECT 23.000 35.900 24.300 36.200 ;
        RECT 24.600 35.900 26.000 36.200 ;
        RECT 27.000 36.200 27.400 36.300 ;
        RECT 27.800 36.200 28.200 39.900 ;
        RECT 27.000 35.900 28.200 36.200 ;
        RECT 24.600 35.800 25.800 35.900 ;
        RECT 18.600 34.900 20.200 35.100 ;
        RECT 16.600 34.800 17.000 34.900 ;
        RECT 16.600 34.200 16.900 34.800 ;
        RECT 10.600 33.600 11.000 33.800 ;
        RECT 10.300 33.100 12.100 33.300 ;
        RECT 12.600 33.100 12.900 33.800 ;
        RECT 10.200 33.000 12.200 33.100 ;
        RECT 10.200 31.100 10.600 33.000 ;
        RECT 11.800 31.100 12.200 33.000 ;
        RECT 12.600 31.100 13.000 33.100 ;
        RECT 15.200 31.100 15.600 33.900 ;
        RECT 16.600 33.800 17.000 34.200 ;
        RECT 16.600 32.800 17.000 33.200 ;
        RECT 17.500 33.100 17.800 34.900 ;
        RECT 19.000 34.800 20.200 34.900 ;
        RECT 20.600 34.800 21.400 35.200 ;
        RECT 18.200 33.800 18.600 34.600 ;
        RECT 22.200 34.200 22.500 35.800 ;
        RECT 24.500 35.200 24.900 35.300 ;
        RECT 25.500 35.200 25.800 35.800 ;
        RECT 24.100 34.900 24.900 35.200 ;
        RECT 24.100 34.800 24.500 34.900 ;
        RECT 25.400 34.800 25.800 35.200 ;
        RECT 24.800 34.300 25.200 34.400 ;
        RECT 23.800 34.200 25.200 34.300 ;
        RECT 21.700 34.100 22.500 34.200 ;
        RECT 21.600 33.900 22.500 34.100 ;
        RECT 23.000 34.000 25.200 34.200 ;
        RECT 25.500 34.200 25.800 34.800 ;
        RECT 23.000 33.900 24.100 34.000 ;
        RECT 25.500 33.900 26.000 34.200 ;
        RECT 16.700 32.400 17.100 32.800 ;
        RECT 17.400 31.100 17.800 33.100 ;
        RECT 21.600 31.100 22.000 33.900 ;
        RECT 23.000 33.800 23.800 33.900 ;
        RECT 23.900 33.400 24.300 33.500 ;
        RECT 23.000 33.100 24.300 33.400 ;
        RECT 24.600 33.200 25.400 33.600 ;
        RECT 23.000 31.100 23.400 33.100 ;
        RECT 25.700 32.900 26.000 33.900 ;
        RECT 26.400 33.800 26.800 34.200 ;
        RECT 27.400 33.800 28.200 34.200 ;
        RECT 26.400 33.600 26.700 33.800 ;
        RECT 26.300 33.200 26.700 33.600 ;
        RECT 27.000 33.400 27.400 33.500 ;
        RECT 27.000 33.100 28.200 33.400 ;
        RECT 29.400 33.100 29.800 39.900 ;
        RECT 25.200 31.100 26.000 32.900 ;
        RECT 27.800 31.100 28.200 33.100 ;
        RECT 28.900 32.800 29.800 33.100 ;
        RECT 28.900 32.200 29.300 32.800 ;
        RECT 28.600 31.800 29.300 32.200 ;
        RECT 28.900 31.100 29.300 31.800 ;
        RECT 31.000 31.100 31.400 39.900 ;
        RECT 32.600 36.200 33.000 39.900 ;
        RECT 34.200 36.400 34.600 39.900 ;
        RECT 32.600 35.900 33.900 36.200 ;
        RECT 34.200 35.900 34.700 36.400 ;
        RECT 33.600 34.900 33.900 35.900 ;
        RECT 33.600 34.500 34.100 34.900 ;
        RECT 33.600 33.700 33.900 34.500 ;
        RECT 34.400 34.200 34.700 35.900 ;
        RECT 34.200 33.800 34.700 34.200 ;
        RECT 32.600 33.400 33.900 33.700 ;
        RECT 31.800 32.400 32.200 33.200 ;
        RECT 32.600 31.100 33.000 33.400 ;
        RECT 34.400 33.100 34.700 33.800 ;
        RECT 36.600 33.100 37.000 39.900 ;
        RECT 38.200 36.200 38.600 39.900 ;
        RECT 39.800 36.400 40.200 39.900 ;
        RECT 41.400 39.600 43.400 39.900 ;
        RECT 38.200 35.900 39.500 36.200 ;
        RECT 39.800 35.900 40.300 36.400 ;
        RECT 41.400 35.900 41.800 39.600 ;
        RECT 42.200 35.900 42.600 39.300 ;
        RECT 43.000 36.200 43.400 39.600 ;
        RECT 44.600 36.200 45.000 39.900 ;
        RECT 43.000 35.900 45.000 36.200 ;
        RECT 39.200 34.900 39.500 35.900 ;
        RECT 39.200 34.500 39.700 34.900 ;
        RECT 37.400 33.400 37.800 34.200 ;
        RECT 39.200 33.700 39.500 34.500 ;
        RECT 40.000 34.200 40.300 35.900 ;
        RECT 42.300 35.600 42.600 35.900 ;
        RECT 39.800 34.100 40.300 34.200 ;
        RECT 41.400 34.800 41.800 35.600 ;
        RECT 42.300 35.300 43.300 35.600 ;
        RECT 43.000 35.200 43.300 35.300 ;
        RECT 44.200 35.200 44.600 35.400 ;
        RECT 43.000 34.800 43.400 35.200 ;
        RECT 44.200 34.900 45.000 35.200 ;
        RECT 44.600 34.800 45.000 34.900 ;
        RECT 41.400 34.100 41.700 34.800 ;
        RECT 39.800 33.800 41.700 34.100 ;
        RECT 38.200 33.400 39.500 33.700 ;
        RECT 34.200 32.800 34.700 33.100 ;
        RECT 36.100 32.800 37.000 33.100 ;
        RECT 34.200 31.100 34.600 32.800 ;
        RECT 36.100 31.100 36.500 32.800 ;
        RECT 38.200 31.100 38.600 33.400 ;
        RECT 40.000 33.100 40.300 33.800 ;
        RECT 43.000 33.100 43.300 34.800 ;
        RECT 46.200 33.100 46.600 39.900 ;
        RECT 50.200 36.400 50.600 39.900 ;
        RECT 50.100 35.900 50.600 36.400 ;
        RECT 51.800 36.200 52.200 39.900 ;
        RECT 50.900 35.900 52.200 36.200 ;
        RECT 52.600 36.200 53.000 39.900 ;
        RECT 54.200 36.400 54.600 39.900 ;
        RECT 52.600 35.900 53.900 36.200 ;
        RECT 54.200 35.900 54.700 36.400 ;
        RECT 55.800 36.200 56.200 39.900 ;
        RECT 57.400 36.400 57.800 39.900 ;
        RECT 59.000 37.500 59.400 39.500 ;
        RECT 61.100 39.200 61.500 39.900 ;
        RECT 61.100 38.800 61.800 39.200 ;
        RECT 55.800 35.900 57.100 36.200 ;
        RECT 57.400 35.900 57.900 36.400 ;
        RECT 50.100 34.200 50.400 35.900 ;
        RECT 50.900 34.900 51.200 35.900 ;
        RECT 50.700 34.500 51.200 34.900 ;
        RECT 47.000 33.400 47.400 34.200 ;
        RECT 47.800 34.100 48.200 34.200 ;
        RECT 50.100 34.100 50.600 34.200 ;
        RECT 47.800 33.800 50.600 34.100 ;
        RECT 39.800 32.800 40.300 33.100 ;
        RECT 39.800 31.100 40.200 32.800 ;
        RECT 42.700 31.100 43.500 33.100 ;
        RECT 45.700 32.800 46.600 33.100 ;
        RECT 50.100 33.100 50.400 33.800 ;
        RECT 50.900 33.700 51.200 34.500 ;
        RECT 53.600 34.900 53.900 35.900 ;
        RECT 53.600 34.500 54.100 34.900 ;
        RECT 53.600 33.700 53.900 34.500 ;
        RECT 54.400 34.200 54.700 35.900 ;
        RECT 56.800 34.900 57.100 35.900 ;
        RECT 56.800 34.500 57.300 34.900 ;
        RECT 54.200 34.100 54.700 34.200 ;
        RECT 55.000 34.100 55.400 34.200 ;
        RECT 54.200 33.800 55.400 34.100 ;
        RECT 50.900 33.400 52.200 33.700 ;
        RECT 50.100 32.800 50.600 33.100 ;
        RECT 45.700 32.200 46.100 32.800 ;
        RECT 45.400 31.800 46.100 32.200 ;
        RECT 45.700 31.100 46.100 31.800 ;
        RECT 50.200 31.100 50.600 32.800 ;
        RECT 51.800 31.100 52.200 33.400 ;
        RECT 52.600 33.400 53.900 33.700 ;
        RECT 52.600 31.100 53.000 33.400 ;
        RECT 54.400 33.100 54.700 33.800 ;
        RECT 56.800 33.700 57.100 34.500 ;
        RECT 57.600 34.200 57.900 35.900 ;
        RECT 59.000 35.800 59.300 37.500 ;
        RECT 61.100 36.400 61.500 38.800 ;
        RECT 65.700 36.400 66.100 39.900 ;
        RECT 67.800 37.500 68.200 39.500 ;
        RECT 61.100 36.100 61.900 36.400 ;
        RECT 59.000 35.500 60.900 35.800 ;
        RECT 59.000 34.400 59.400 35.200 ;
        RECT 59.800 34.400 60.200 35.200 ;
        RECT 60.600 34.500 60.900 35.500 ;
        RECT 57.400 33.800 57.900 34.200 ;
        RECT 60.600 34.100 61.300 34.500 ;
        RECT 61.600 34.200 61.900 36.100 ;
        RECT 65.300 36.100 66.100 36.400 ;
        RECT 62.200 35.100 62.600 35.600 ;
        RECT 62.200 34.800 63.300 35.100 ;
        RECT 60.600 33.900 61.100 34.100 ;
        RECT 54.200 32.800 54.700 33.100 ;
        RECT 55.800 33.400 57.100 33.700 ;
        RECT 54.200 31.100 54.600 32.800 ;
        RECT 55.800 31.100 56.200 33.400 ;
        RECT 57.600 33.100 57.900 33.800 ;
        RECT 57.400 32.800 57.900 33.100 ;
        RECT 59.000 33.600 61.100 33.900 ;
        RECT 61.600 33.800 62.600 34.200 ;
        RECT 63.000 34.100 63.300 34.800 ;
        RECT 65.300 34.200 65.600 36.100 ;
        RECT 67.900 35.800 68.200 37.500 ;
        RECT 69.900 36.200 70.300 39.900 ;
        RECT 70.600 36.800 71.000 37.200 ;
        RECT 70.700 36.200 71.000 36.800 ;
        RECT 71.800 36.200 72.200 39.900 ;
        RECT 73.400 36.200 73.800 39.900 ;
        RECT 69.900 35.900 70.400 36.200 ;
        RECT 70.700 35.900 71.400 36.200 ;
        RECT 71.800 35.900 73.800 36.200 ;
        RECT 74.200 35.900 74.600 39.900 ;
        RECT 76.300 39.200 76.700 39.900 ;
        RECT 75.800 38.800 76.700 39.200 ;
        RECT 76.300 36.200 76.700 38.800 ;
        RECT 77.000 36.800 77.800 37.200 ;
        RECT 78.600 36.800 79.000 37.200 ;
        RECT 77.100 36.200 77.400 36.800 ;
        RECT 78.600 36.200 78.900 36.800 ;
        RECT 79.300 36.200 79.700 39.900 ;
        RECT 76.300 35.900 76.800 36.200 ;
        RECT 77.100 36.100 77.800 36.200 ;
        RECT 78.200 36.100 78.900 36.200 ;
        RECT 77.100 35.900 78.900 36.100 ;
        RECT 79.200 35.900 79.700 36.200 ;
        RECT 82.700 36.200 83.100 39.900 ;
        RECT 83.400 36.800 83.800 37.200 ;
        RECT 83.500 36.200 83.800 36.800 ;
        RECT 82.700 35.900 83.200 36.200 ;
        RECT 83.500 35.900 84.200 36.200 ;
        RECT 66.300 35.500 68.200 35.800 ;
        RECT 66.300 34.500 66.600 35.500 ;
        RECT 70.100 35.200 70.400 35.900 ;
        RECT 71.000 35.800 71.400 35.900 ;
        RECT 72.200 35.200 72.600 35.400 ;
        RECT 74.200 35.200 74.500 35.900 ;
        RECT 64.600 34.100 65.600 34.200 ;
        RECT 65.900 34.100 66.600 34.500 ;
        RECT 67.800 35.100 68.200 35.200 ;
        RECT 68.600 35.100 69.000 35.200 ;
        RECT 67.800 34.800 69.000 35.100 ;
        RECT 67.800 34.400 68.200 34.800 ;
        RECT 69.400 34.400 69.800 35.200 ;
        RECT 70.100 34.800 70.600 35.200 ;
        RECT 71.800 34.900 72.600 35.200 ;
        RECT 73.400 34.900 74.600 35.200 ;
        RECT 71.800 34.800 72.200 34.900 ;
        RECT 70.100 34.200 70.400 34.800 ;
        RECT 63.000 33.800 65.600 34.100 ;
        RECT 57.400 31.100 57.800 32.800 ;
        RECT 59.000 32.500 59.300 33.600 ;
        RECT 61.600 33.500 61.900 33.800 ;
        RECT 61.500 33.300 61.900 33.500 ;
        RECT 61.100 33.000 61.900 33.300 ;
        RECT 65.300 33.500 65.600 33.800 ;
        RECT 66.100 33.900 66.600 34.100 ;
        RECT 68.600 34.100 69.000 34.200 ;
        RECT 66.100 33.600 68.200 33.900 ;
        RECT 68.600 33.800 69.400 34.100 ;
        RECT 70.100 33.800 71.400 34.200 ;
        RECT 71.800 34.100 72.200 34.200 ;
        RECT 72.600 34.100 73.000 34.600 ;
        RECT 71.800 33.800 73.000 34.100 ;
        RECT 69.000 33.600 69.400 33.800 ;
        RECT 65.300 33.300 65.700 33.500 ;
        RECT 65.300 33.200 66.100 33.300 ;
        RECT 65.300 33.000 66.600 33.200 ;
        RECT 59.000 31.500 59.400 32.500 ;
        RECT 61.100 31.500 61.500 33.000 ;
        RECT 65.700 32.800 66.600 33.000 ;
        RECT 65.700 31.500 66.100 32.800 ;
        RECT 67.900 32.500 68.200 33.600 ;
        RECT 68.700 33.100 70.500 33.300 ;
        RECT 71.000 33.100 71.300 33.800 ;
        RECT 73.400 33.100 73.700 34.900 ;
        RECT 74.200 34.800 74.600 34.900 ;
        RECT 75.800 34.400 76.200 35.200 ;
        RECT 76.500 34.200 76.800 35.900 ;
        RECT 77.400 35.800 78.600 35.900 ;
        RECT 79.200 34.200 79.500 35.900 ;
        RECT 79.800 34.400 80.200 35.200 ;
        RECT 82.200 34.400 82.600 35.200 ;
        RECT 82.900 34.200 83.200 35.900 ;
        RECT 83.800 35.800 84.200 35.900 ;
        RECT 84.600 35.800 85.000 36.600 ;
        RECT 83.800 35.200 84.100 35.800 ;
        RECT 83.800 34.800 84.200 35.200 ;
        RECT 75.000 34.100 75.400 34.200 ;
        RECT 75.000 33.800 75.800 34.100 ;
        RECT 76.500 33.800 77.800 34.200 ;
        RECT 78.200 33.800 79.500 34.200 ;
        RECT 80.600 34.100 81.000 34.200 ;
        RECT 80.200 33.800 81.000 34.100 ;
        RECT 81.400 34.100 81.800 34.200 ;
        RECT 81.400 33.800 82.200 34.100 ;
        RECT 82.900 33.800 84.200 34.200 ;
        RECT 75.400 33.600 75.800 33.800 ;
        RECT 67.800 31.500 68.200 32.500 ;
        RECT 68.600 33.000 70.600 33.100 ;
        RECT 68.600 31.100 69.000 33.000 ;
        RECT 70.200 31.100 70.600 33.000 ;
        RECT 71.000 31.100 71.400 33.100 ;
        RECT 73.400 31.100 73.800 33.100 ;
        RECT 74.200 32.800 74.600 33.200 ;
        RECT 75.100 33.100 76.900 33.300 ;
        RECT 77.400 33.100 77.700 33.800 ;
        RECT 78.300 33.100 78.600 33.800 ;
        RECT 80.200 33.600 80.600 33.800 ;
        RECT 81.800 33.600 82.200 33.800 ;
        RECT 79.100 33.100 80.900 33.300 ;
        RECT 81.500 33.100 83.300 33.300 ;
        RECT 83.800 33.200 84.100 33.800 ;
        RECT 75.000 33.000 77.000 33.100 ;
        RECT 74.100 32.400 74.500 32.800 ;
        RECT 75.000 31.100 75.400 33.000 ;
        RECT 76.600 31.100 77.000 33.000 ;
        RECT 77.400 31.100 77.800 33.100 ;
        RECT 78.200 31.100 78.600 33.100 ;
        RECT 79.000 33.000 81.000 33.100 ;
        RECT 79.000 31.100 79.400 33.000 ;
        RECT 80.600 31.100 81.000 33.000 ;
        RECT 81.400 33.000 83.400 33.100 ;
        RECT 81.400 31.100 81.800 33.000 ;
        RECT 83.000 31.100 83.400 33.000 ;
        RECT 83.800 31.100 84.200 33.200 ;
        RECT 85.400 33.100 85.800 39.900 ;
        RECT 88.300 37.200 88.700 39.900 ;
        RECT 88.300 36.800 89.000 37.200 ;
        RECT 88.300 36.300 88.700 36.800 ;
        RECT 87.800 35.900 88.700 36.300 ;
        RECT 89.400 35.900 89.800 39.900 ;
        RECT 90.200 36.200 90.600 39.900 ;
        RECT 91.800 36.200 92.200 39.900 ;
        RECT 90.200 35.900 92.200 36.200 ;
        RECT 92.900 36.300 93.300 39.900 ;
        RECT 92.900 35.900 93.800 36.300 ;
        RECT 96.300 36.200 96.700 39.900 ;
        RECT 97.000 36.800 97.400 37.200 ;
        RECT 97.100 36.200 97.400 36.800 ;
        RECT 96.300 35.900 96.800 36.200 ;
        RECT 97.100 35.900 97.800 36.200 ;
        RECT 98.200 35.900 98.600 39.900 ;
        RECT 99.000 36.200 99.400 39.900 ;
        RECT 100.600 36.200 101.000 39.900 ;
        RECT 99.000 35.900 101.000 36.200 ;
        RECT 87.900 34.200 88.200 35.900 ;
        RECT 88.600 34.800 89.000 35.600 ;
        RECT 89.500 35.200 89.800 35.900 ;
        RECT 91.400 35.200 91.800 35.400 ;
        RECT 89.400 34.900 90.600 35.200 ;
        RECT 91.400 34.900 92.200 35.200 ;
        RECT 89.400 34.800 89.800 34.900 ;
        RECT 90.200 34.800 90.600 34.900 ;
        RECT 91.800 34.800 92.200 34.900 ;
        RECT 92.600 34.800 93.000 35.600 ;
        RECT 93.400 35.100 93.700 35.900 ;
        RECT 93.400 34.800 95.300 35.100 ;
        RECT 86.200 33.400 86.600 34.200 ;
        RECT 87.800 33.800 88.200 34.200 ;
        RECT 84.900 32.800 85.800 33.100 ;
        RECT 84.900 31.100 85.300 32.800 ;
        RECT 87.000 32.400 87.400 33.200 ;
        RECT 87.900 32.100 88.200 33.800 ;
        RECT 89.400 32.800 89.800 33.200 ;
        RECT 90.300 33.100 90.600 34.800 ;
        RECT 91.000 33.800 91.400 34.600 ;
        RECT 93.400 34.200 93.700 34.800 ;
        RECT 95.000 34.200 95.300 34.800 ;
        RECT 95.800 34.400 96.200 35.200 ;
        RECT 96.500 34.200 96.800 35.900 ;
        RECT 97.400 35.800 97.800 35.900 ;
        RECT 98.300 35.200 98.600 35.900 ;
        RECT 103.000 35.800 103.400 36.600 ;
        RECT 103.800 36.100 104.200 39.900 ;
        RECT 104.600 36.800 105.000 37.200 ;
        RECT 104.600 36.100 104.900 36.800 ;
        RECT 103.800 35.800 104.900 36.100 ;
        RECT 100.200 35.200 100.600 35.400 ;
        RECT 98.200 34.900 99.400 35.200 ;
        RECT 100.200 35.100 101.000 35.200 ;
        RECT 101.400 35.100 101.800 35.200 ;
        RECT 100.200 34.900 101.800 35.100 ;
        RECT 98.200 34.800 98.600 34.900 ;
        RECT 93.400 33.800 93.800 34.200 ;
        RECT 95.000 34.100 95.400 34.200 ;
        RECT 95.000 33.800 95.800 34.100 ;
        RECT 96.500 33.800 97.800 34.200 ;
        RECT 89.500 32.400 89.900 32.800 ;
        RECT 87.800 31.100 88.200 32.100 ;
        RECT 90.200 31.100 90.600 33.100 ;
        RECT 93.400 32.100 93.700 33.800 ;
        RECT 95.400 33.600 95.800 33.800 ;
        RECT 94.200 32.400 94.600 33.200 ;
        RECT 95.100 33.100 96.900 33.300 ;
        RECT 97.400 33.100 97.700 33.800 ;
        RECT 95.000 33.000 97.000 33.100 ;
        RECT 93.400 31.100 93.800 32.100 ;
        RECT 95.000 31.100 95.400 33.000 ;
        RECT 96.600 31.100 97.000 33.000 ;
        RECT 97.400 31.100 97.800 33.100 ;
        RECT 98.200 32.800 98.600 33.200 ;
        RECT 99.100 33.100 99.400 34.900 ;
        RECT 100.600 34.800 101.800 34.900 ;
        RECT 99.800 34.100 100.200 34.600 ;
        RECT 102.200 34.100 102.600 34.200 ;
        RECT 99.800 33.800 102.600 34.100 ;
        RECT 103.800 33.100 104.200 35.800 ;
        RECT 104.600 33.400 105.000 34.200 ;
        RECT 98.300 32.400 98.700 32.800 ;
        RECT 99.000 31.100 99.400 33.100 ;
        RECT 103.300 32.800 104.200 33.100 ;
        RECT 103.300 31.100 103.700 32.800 ;
        RECT 105.400 31.100 105.800 39.900 ;
        RECT 108.100 38.200 108.500 39.900 ;
        RECT 108.100 37.800 109.000 38.200 ;
        RECT 107.400 36.800 107.800 37.200 ;
        RECT 107.400 36.200 107.700 36.800 ;
        RECT 108.100 36.200 108.500 37.800 ;
        RECT 107.000 35.900 107.700 36.200 ;
        RECT 108.000 35.900 108.500 36.200 ;
        RECT 110.500 36.300 110.900 39.900 ;
        RECT 113.400 37.900 113.800 39.900 ;
        RECT 110.500 35.900 111.400 36.300 ;
        RECT 107.000 35.800 107.400 35.900 ;
        RECT 108.000 34.200 108.300 35.900 ;
        RECT 108.600 35.100 109.000 35.200 ;
        RECT 109.400 35.100 109.800 35.200 ;
        RECT 108.600 34.800 109.800 35.100 ;
        RECT 110.200 34.800 110.600 35.600 ;
        RECT 111.000 35.100 111.300 35.900 ;
        RECT 113.500 35.800 113.800 37.900 ;
        RECT 115.000 35.900 115.400 39.900 ;
        RECT 117.100 36.200 117.500 39.900 ;
        RECT 117.800 36.800 118.200 37.200 ;
        RECT 117.900 36.200 118.200 36.800 ;
        RECT 117.100 35.900 117.600 36.200 ;
        RECT 117.900 35.900 118.600 36.200 ;
        RECT 113.500 35.500 114.700 35.800 ;
        RECT 111.000 34.800 112.100 35.100 ;
        RECT 113.400 34.800 113.800 35.200 ;
        RECT 108.600 34.400 109.000 34.800 ;
        RECT 111.000 34.200 111.300 34.800 ;
        RECT 111.800 34.200 112.100 34.800 ;
        RECT 106.200 33.400 106.600 34.200 ;
        RECT 107.000 33.800 108.300 34.200 ;
        RECT 109.400 34.100 109.800 34.200 ;
        RECT 109.000 33.800 109.800 34.100 ;
        RECT 111.000 33.800 111.400 34.200 ;
        RECT 111.800 33.800 112.200 34.200 ;
        RECT 112.600 33.800 113.000 34.600 ;
        RECT 113.500 34.400 113.800 34.800 ;
        RECT 113.500 34.100 114.000 34.400 ;
        RECT 113.600 34.000 114.000 34.100 ;
        RECT 114.400 33.800 114.700 35.500 ;
        RECT 115.100 35.200 115.400 35.900 ;
        RECT 115.000 34.800 115.400 35.200 ;
        RECT 115.800 35.100 116.200 35.200 ;
        RECT 116.600 35.100 117.000 35.200 ;
        RECT 115.800 34.800 117.000 35.100 ;
        RECT 107.100 33.100 107.400 33.800 ;
        RECT 109.000 33.600 109.400 33.800 ;
        RECT 107.900 33.100 109.700 33.300 ;
        RECT 107.000 31.100 107.400 33.100 ;
        RECT 107.800 33.000 109.800 33.100 ;
        RECT 107.800 31.100 108.200 33.000 ;
        RECT 109.400 31.100 109.800 33.000 ;
        RECT 111.000 32.100 111.300 33.800 ;
        RECT 114.400 33.700 114.800 33.800 ;
        RECT 113.300 33.500 114.800 33.700 ;
        RECT 112.700 33.400 114.800 33.500 ;
        RECT 112.700 33.200 113.600 33.400 ;
        RECT 111.800 32.400 112.200 33.200 ;
        RECT 112.700 33.100 113.000 33.200 ;
        RECT 115.100 33.100 115.400 34.800 ;
        RECT 116.600 34.400 117.000 34.800 ;
        RECT 117.300 34.200 117.600 35.900 ;
        RECT 118.200 35.800 118.600 35.900 ;
        RECT 119.000 35.100 119.400 35.200 ;
        RECT 119.800 35.100 120.200 39.900 ;
        RECT 120.600 35.800 121.000 36.600 ;
        RECT 121.400 35.600 121.800 39.900 ;
        RECT 123.500 36.200 123.900 39.900 ;
        RECT 124.600 36.200 125.000 39.900 ;
        RECT 126.200 36.200 126.600 39.900 ;
        RECT 123.500 35.900 124.200 36.200 ;
        RECT 124.600 35.900 126.600 36.200 ;
        RECT 127.000 35.900 127.400 39.900 ;
        RECT 129.100 39.200 129.500 39.900 ;
        RECT 128.600 38.800 129.500 39.200 ;
        RECT 129.100 36.300 129.500 38.800 ;
        RECT 128.600 35.900 129.500 36.300 ;
        RECT 130.500 36.200 130.900 39.900 ;
        RECT 130.200 35.900 130.900 36.200 ;
        RECT 121.400 35.400 123.400 35.600 ;
        RECT 121.400 35.300 123.500 35.400 ;
        RECT 119.000 34.800 120.200 35.100 ;
        RECT 123.100 35.000 123.500 35.300 ;
        RECT 123.900 35.200 124.200 35.900 ;
        RECT 125.000 35.200 125.400 35.400 ;
        RECT 127.000 35.200 127.300 35.900 ;
        RECT 115.800 34.100 116.200 34.200 ;
        RECT 115.800 33.800 116.600 34.100 ;
        RECT 117.300 33.800 118.600 34.200 ;
        RECT 116.200 33.600 116.600 33.800 ;
        RECT 115.900 33.100 117.700 33.300 ;
        RECT 118.200 33.100 118.500 33.800 ;
        RECT 119.000 33.400 119.400 34.200 ;
        RECT 119.800 33.100 120.200 34.800 ;
        RECT 122.400 34.200 122.800 34.600 ;
        RECT 122.200 33.800 122.700 34.200 ;
        RECT 123.200 33.500 123.500 35.000 ;
        RECT 123.800 34.800 124.200 35.200 ;
        RECT 124.600 34.900 125.400 35.200 ;
        RECT 126.200 34.900 127.400 35.200 ;
        RECT 124.600 34.800 125.000 34.900 ;
        RECT 123.900 34.100 124.200 34.800 ;
        RECT 125.400 34.100 125.800 34.600 ;
        RECT 123.800 33.800 125.800 34.100 ;
        RECT 126.200 34.100 126.500 34.900 ;
        RECT 127.000 34.800 127.400 34.900 ;
        RECT 128.700 34.200 129.000 35.900 ;
        RECT 129.400 35.100 129.800 35.600 ;
        RECT 130.200 35.200 130.500 35.900 ;
        RECT 132.600 35.600 133.000 39.900 ;
        RECT 131.000 35.400 133.000 35.600 ;
        RECT 130.900 35.300 133.000 35.400 ;
        RECT 130.200 35.100 130.600 35.200 ;
        RECT 129.400 34.800 130.600 35.100 ;
        RECT 130.900 35.000 131.300 35.300 ;
        RECT 126.200 33.800 128.100 34.100 ;
        RECT 128.600 33.800 129.000 34.200 ;
        RECT 122.300 33.200 123.500 33.500 ;
        RECT 111.000 31.100 111.400 32.100 ;
        RECT 112.600 31.100 113.000 33.100 ;
        RECT 114.700 32.600 115.400 33.100 ;
        RECT 115.800 33.000 117.800 33.100 ;
        RECT 114.700 32.200 115.100 32.600 ;
        RECT 114.700 31.800 115.400 32.200 ;
        RECT 114.700 31.100 115.100 31.800 ;
        RECT 115.800 31.100 116.200 33.000 ;
        RECT 117.400 31.100 117.800 33.000 ;
        RECT 118.200 31.100 118.600 33.100 ;
        RECT 119.800 32.800 120.700 33.100 ;
        RECT 120.300 31.100 120.700 32.800 ;
        RECT 121.400 32.400 121.800 33.200 ;
        RECT 122.300 32.100 122.600 33.200 ;
        RECT 123.900 33.100 124.200 33.800 ;
        RECT 122.200 31.100 122.600 32.100 ;
        RECT 123.800 31.100 124.200 33.100 ;
        RECT 126.200 33.100 126.500 33.800 ;
        RECT 127.800 33.200 128.100 33.800 ;
        RECT 126.200 31.100 126.600 33.100 ;
        RECT 127.000 32.800 127.400 33.200 ;
        RECT 126.900 32.400 127.300 32.800 ;
        RECT 127.800 32.400 128.200 33.200 ;
        RECT 128.700 32.100 129.000 33.800 ;
        RECT 128.600 31.100 129.000 32.100 ;
        RECT 130.200 33.100 130.500 34.800 ;
        RECT 130.900 33.500 131.200 35.000 ;
        RECT 131.600 34.200 132.000 34.600 ;
        RECT 131.700 33.800 132.200 34.200 ;
        RECT 130.900 33.200 132.100 33.500 ;
        RECT 130.200 31.100 130.600 33.100 ;
        RECT 131.800 32.100 132.100 33.200 ;
        RECT 132.600 32.400 133.000 33.200 ;
        RECT 131.800 31.100 132.200 32.100 ;
        RECT 133.400 31.100 133.800 39.900 ;
        RECT 135.000 37.900 135.400 39.900 ;
        RECT 135.100 37.800 135.400 37.900 ;
        RECT 136.600 37.900 137.000 39.900 ;
        RECT 136.600 37.800 136.900 37.900 ;
        RECT 135.100 37.500 136.900 37.800 ;
        RECT 135.100 36.200 135.400 37.500 ;
        RECT 135.800 36.400 136.200 37.200 ;
        RECT 138.500 36.200 138.900 39.900 ;
        RECT 135.000 35.800 135.400 36.200 ;
        RECT 135.100 34.200 135.400 35.800 ;
        RECT 137.400 35.400 137.800 36.200 ;
        RECT 138.200 35.900 138.900 36.200 ;
        RECT 138.200 35.200 138.500 35.900 ;
        RECT 140.600 35.600 141.000 39.900 ;
        RECT 141.700 39.200 142.100 39.900 ;
        RECT 141.400 38.800 142.100 39.200 ;
        RECT 141.700 36.300 142.100 38.800 ;
        RECT 141.700 35.900 142.600 36.300 ;
        RECT 139.000 35.400 141.000 35.600 ;
        RECT 138.900 35.300 141.000 35.400 ;
        RECT 136.200 34.800 137.000 35.200 ;
        RECT 138.200 34.800 138.600 35.200 ;
        RECT 138.900 35.000 139.300 35.300 ;
        RECT 134.200 33.400 134.600 34.200 ;
        RECT 135.100 34.100 135.900 34.200 ;
        RECT 135.100 33.900 136.000 34.100 ;
        RECT 135.600 31.100 136.000 33.900 ;
        RECT 138.200 33.100 138.500 34.800 ;
        RECT 138.900 33.500 139.200 35.000 ;
        RECT 141.400 34.800 141.800 35.600 ;
        RECT 139.600 34.200 140.000 34.600 ;
        RECT 142.200 34.200 142.500 35.900 ;
        RECT 143.800 35.100 144.200 35.200 ;
        RECT 144.600 35.100 145.000 39.900 ;
        RECT 146.500 36.200 146.900 39.900 ;
        RECT 143.800 34.800 145.000 35.100 ;
        RECT 139.700 33.800 140.200 34.200 ;
        RECT 142.200 33.800 142.600 34.200 ;
        RECT 138.900 33.200 140.100 33.500 ;
        RECT 138.200 31.100 138.600 33.100 ;
        RECT 139.800 32.100 140.100 33.200 ;
        RECT 140.600 33.100 141.000 33.200 ;
        RECT 141.400 33.100 141.800 33.200 ;
        RECT 140.600 32.800 141.800 33.100 ;
        RECT 140.600 32.400 141.000 32.800 ;
        RECT 142.200 32.100 142.500 33.800 ;
        RECT 144.600 33.100 145.000 34.800 ;
        RECT 144.100 32.800 145.000 33.100 ;
        RECT 146.200 35.900 146.900 36.200 ;
        RECT 146.200 35.200 146.500 35.900 ;
        RECT 148.600 35.600 149.000 39.900 ;
        RECT 147.000 35.400 149.000 35.600 ;
        RECT 146.900 35.300 149.000 35.400 ;
        RECT 146.200 34.800 146.600 35.200 ;
        RECT 146.900 35.000 147.300 35.300 ;
        RECT 146.200 33.100 146.500 34.800 ;
        RECT 146.900 33.500 147.200 35.000 ;
        RECT 146.900 33.200 148.100 33.500 ;
        RECT 139.800 31.100 140.200 32.100 ;
        RECT 142.200 31.100 142.600 32.100 ;
        RECT 144.100 31.100 144.500 32.800 ;
        RECT 146.200 31.100 146.600 33.100 ;
        RECT 147.800 32.100 148.100 33.200 ;
        RECT 147.800 31.100 148.200 32.100 ;
        RECT 0.600 27.900 1.000 29.900 ;
        RECT 2.800 28.100 3.600 29.900 ;
        RECT 0.600 27.600 1.800 27.900 ;
        RECT 1.400 27.500 1.800 27.600 ;
        RECT 2.100 27.400 2.500 27.800 ;
        RECT 2.100 27.200 2.400 27.400 ;
        RECT 0.600 26.800 1.400 27.200 ;
        RECT 2.000 26.800 2.400 27.200 ;
        RECT 2.800 26.400 3.100 28.100 ;
        RECT 5.400 27.900 5.800 29.900 ;
        RECT 3.400 27.700 4.200 27.800 ;
        RECT 3.400 27.400 4.400 27.700 ;
        RECT 4.700 27.600 5.800 27.900 ;
        RECT 6.800 29.200 7.200 29.900 ;
        RECT 6.800 28.800 7.400 29.200 ;
        RECT 4.700 27.500 5.100 27.600 ;
        RECT 4.100 27.200 4.400 27.400 ;
        RECT 3.400 26.700 3.800 27.100 ;
        RECT 4.100 26.900 5.800 27.200 ;
        RECT 6.800 27.100 7.200 28.800 ;
        RECT 11.000 27.900 11.400 29.900 ;
        RECT 11.700 28.200 12.100 28.600 ;
        RECT 11.800 28.100 12.200 28.200 ;
        RECT 12.600 28.100 13.000 28.600 ;
        RECT 5.000 26.800 5.800 26.900 ;
        RECT 6.300 26.900 7.200 27.100 ;
        RECT 6.300 26.800 7.100 26.900 ;
        RECT 2.600 26.200 3.100 26.400 ;
        RECT 2.200 26.100 3.100 26.200 ;
        RECT 3.500 26.400 3.800 26.700 ;
        RECT 3.500 26.100 4.800 26.400 ;
        RECT 2.200 25.800 2.900 26.100 ;
        RECT 4.400 26.000 4.800 26.100 ;
        RECT 2.600 25.100 2.900 25.800 ;
        RECT 3.300 25.700 3.700 25.800 ;
        RECT 3.300 25.400 5.000 25.700 ;
        RECT 4.700 25.100 5.000 25.400 ;
        RECT 6.300 25.200 6.600 26.800 ;
        RECT 10.200 26.400 10.600 27.200 ;
        RECT 7.400 25.800 8.200 26.200 ;
        RECT 9.400 26.100 9.800 26.200 ;
        RECT 11.000 26.100 11.300 27.900 ;
        RECT 11.800 27.800 13.000 28.100 ;
        RECT 13.400 28.100 13.800 29.900 ;
        RECT 14.300 28.200 14.700 28.600 ;
        RECT 14.200 28.100 14.600 28.200 ;
        RECT 13.400 27.800 14.600 28.100 ;
        RECT 15.000 27.900 15.400 29.900 ;
        RECT 19.200 29.200 19.600 29.900 ;
        RECT 19.000 28.800 19.600 29.200 ;
        RECT 13.400 27.100 13.800 27.800 ;
        RECT 14.200 27.100 14.600 27.200 ;
        RECT 13.400 26.800 14.600 27.100 ;
        RECT 11.800 26.100 12.200 26.200 ;
        RECT 9.400 25.800 10.200 26.100 ;
        RECT 11.000 25.800 12.200 26.100 ;
        RECT 9.800 25.600 10.200 25.800 ;
        RECT 0.600 24.800 1.800 25.100 ;
        RECT 2.600 24.800 3.600 25.100 ;
        RECT 0.600 21.100 1.000 24.800 ;
        RECT 1.400 24.700 1.800 24.800 ;
        RECT 2.800 24.200 3.600 24.800 ;
        RECT 4.700 24.800 5.800 25.100 ;
        RECT 6.200 24.800 6.600 25.200 ;
        RECT 8.600 24.800 9.000 25.600 ;
        RECT 11.800 25.100 12.100 25.800 ;
        RECT 9.400 24.800 11.400 25.100 ;
        RECT 4.700 24.700 5.100 24.800 ;
        RECT 2.800 23.800 4.200 24.200 ;
        RECT 2.800 21.100 3.600 23.800 ;
        RECT 5.400 21.100 5.800 24.800 ;
        RECT 6.300 23.500 6.600 24.800 ;
        RECT 7.000 24.100 7.400 24.600 ;
        RECT 8.600 24.100 9.000 24.200 ;
        RECT 7.000 23.800 9.000 24.100 ;
        RECT 6.300 23.200 8.100 23.500 ;
        RECT 6.300 23.100 6.600 23.200 ;
        RECT 6.200 21.100 6.600 23.100 ;
        RECT 7.800 23.100 8.100 23.200 ;
        RECT 7.800 21.100 8.200 23.100 ;
        RECT 9.400 21.100 9.800 24.800 ;
        RECT 11.000 21.100 11.400 24.800 ;
        RECT 11.800 21.100 12.200 25.100 ;
        RECT 13.400 21.100 13.800 26.800 ;
        RECT 14.200 26.100 14.600 26.200 ;
        RECT 15.100 26.100 15.400 27.900 ;
        RECT 15.800 26.400 16.200 27.200 ;
        RECT 19.200 27.100 19.600 28.800 ;
        RECT 21.900 28.200 22.300 29.900 ;
        RECT 21.400 27.900 22.300 28.200 ;
        RECT 21.400 27.100 21.800 27.900 ;
        RECT 22.200 27.100 22.600 27.200 ;
        RECT 23.600 27.100 24.000 29.900 ;
        RECT 26.800 27.100 27.200 29.900 ;
        RECT 30.200 28.200 30.600 29.900 ;
        RECT 30.100 27.900 30.600 28.200 ;
        RECT 30.100 27.200 30.400 27.900 ;
        RECT 31.800 27.600 32.200 29.900 ;
        RECT 30.900 27.300 32.200 27.600 ;
        RECT 32.600 27.600 33.000 29.900 ;
        RECT 34.200 28.200 34.600 29.900 ;
        RECT 35.800 29.600 37.800 29.900 ;
        RECT 34.200 27.900 34.700 28.200 ;
        RECT 35.800 27.900 36.200 29.600 ;
        RECT 36.600 27.900 37.000 29.300 ;
        RECT 37.400 28.000 37.800 29.600 ;
        RECT 39.000 28.000 39.400 29.900 ;
        RECT 37.400 27.900 39.400 28.000 ;
        RECT 32.600 27.300 33.900 27.600 ;
        RECT 19.200 26.900 20.100 27.100 ;
        RECT 19.300 26.800 20.100 26.900 ;
        RECT 16.600 26.100 17.000 26.200 ;
        RECT 14.200 25.800 15.400 26.100 ;
        RECT 16.200 25.800 17.000 26.100 ;
        RECT 18.200 25.800 19.000 26.200 ;
        RECT 14.300 25.100 14.600 25.800 ;
        RECT 16.200 25.600 16.600 25.800 ;
        RECT 14.200 21.100 14.600 25.100 ;
        RECT 15.000 24.800 17.000 25.100 ;
        RECT 17.400 24.800 17.800 25.600 ;
        RECT 19.800 25.200 20.100 26.800 ;
        RECT 21.400 26.800 22.600 27.100 ;
        RECT 23.100 26.900 24.000 27.100 ;
        RECT 26.300 26.900 27.200 27.100 ;
        RECT 29.400 27.100 29.800 27.200 ;
        RECT 30.100 27.100 30.600 27.200 ;
        RECT 23.100 26.800 23.900 26.900 ;
        RECT 26.300 26.800 27.100 26.900 ;
        RECT 29.400 26.800 30.600 27.100 ;
        RECT 19.800 24.800 20.200 25.200 ;
        RECT 15.000 21.100 15.400 24.800 ;
        RECT 16.600 21.100 17.000 24.800 ;
        RECT 19.000 23.800 19.400 24.600 ;
        RECT 19.800 23.500 20.100 24.800 ;
        RECT 18.300 23.200 20.100 23.500 ;
        RECT 18.300 23.100 18.600 23.200 ;
        RECT 18.200 21.100 18.600 23.100 ;
        RECT 19.800 23.100 20.100 23.200 ;
        RECT 19.800 21.100 20.200 23.100 ;
        RECT 21.400 21.100 21.800 26.800 ;
        RECT 23.100 25.200 23.400 26.800 ;
        RECT 26.300 25.200 26.600 26.800 ;
        RECT 23.000 24.800 23.400 25.200 ;
        RECT 26.200 24.800 26.600 25.200 ;
        RECT 23.100 23.500 23.400 24.800 ;
        RECT 23.800 23.800 24.200 24.600 ;
        RECT 26.300 23.500 26.600 24.800 ;
        RECT 30.100 25.100 30.400 26.800 ;
        RECT 30.900 26.500 31.200 27.300 ;
        RECT 30.700 26.100 31.200 26.500 ;
        RECT 30.900 25.100 31.200 26.100 ;
        RECT 33.600 26.500 33.900 27.300 ;
        RECT 34.400 27.200 34.700 27.900 ;
        RECT 36.600 27.200 36.900 27.900 ;
        RECT 37.500 27.700 39.300 27.900 ;
        RECT 38.600 27.200 39.000 27.400 ;
        RECT 34.200 26.800 34.700 27.200 ;
        RECT 35.000 27.100 35.400 27.200 ;
        RECT 35.800 27.100 36.200 27.200 ;
        RECT 35.000 26.800 36.200 27.100 ;
        RECT 36.600 26.900 37.800 27.200 ;
        RECT 38.600 26.900 39.400 27.200 ;
        RECT 40.400 27.100 40.800 29.900 ;
        RECT 37.400 26.800 37.800 26.900 ;
        RECT 39.000 26.800 39.400 26.900 ;
        RECT 39.900 26.900 40.800 27.100 ;
        RECT 44.800 27.100 45.200 29.900 ;
        RECT 47.000 28.200 47.400 29.900 ;
        RECT 46.900 27.900 47.400 28.200 ;
        RECT 46.900 27.200 47.200 27.900 ;
        RECT 48.600 27.600 49.000 29.900 ;
        RECT 47.700 27.300 49.000 27.600 ;
        RECT 46.200 27.100 46.600 27.200 ;
        RECT 46.900 27.100 47.400 27.200 ;
        RECT 44.800 26.900 45.700 27.100 ;
        RECT 39.900 26.800 40.700 26.900 ;
        RECT 44.900 26.800 45.700 26.900 ;
        RECT 46.200 26.800 47.400 27.100 ;
        RECT 33.600 26.100 34.100 26.500 ;
        RECT 33.600 25.100 33.900 26.100 ;
        RECT 34.400 25.200 34.700 26.800 ;
        RECT 35.800 26.400 36.200 26.800 ;
        RECT 36.600 25.800 37.000 26.600 ;
        RECT 30.100 24.600 30.600 25.100 ;
        RECT 30.900 24.800 32.200 25.100 ;
        RECT 27.000 23.800 27.400 24.600 ;
        RECT 23.100 23.200 24.900 23.500 ;
        RECT 23.100 23.100 23.400 23.200 ;
        RECT 23.000 21.100 23.400 23.100 ;
        RECT 24.600 23.100 24.900 23.200 ;
        RECT 26.300 23.200 28.100 23.500 ;
        RECT 26.300 23.100 26.600 23.200 ;
        RECT 24.600 21.100 25.000 23.100 ;
        RECT 26.200 21.100 26.600 23.100 ;
        RECT 27.800 23.100 28.100 23.200 ;
        RECT 27.800 21.100 28.200 23.100 ;
        RECT 30.200 21.100 30.600 24.600 ;
        RECT 31.800 21.100 32.200 24.800 ;
        RECT 32.600 24.800 33.900 25.100 ;
        RECT 32.600 21.100 33.000 24.800 ;
        RECT 34.200 24.600 34.700 25.200 ;
        RECT 37.500 25.100 37.800 26.800 ;
        RECT 38.200 25.800 38.600 26.600 ;
        RECT 39.900 25.200 40.200 26.800 ;
        RECT 34.200 21.100 34.600 24.600 ;
        RECT 37.100 22.200 38.100 25.100 ;
        RECT 39.800 24.800 40.200 25.200 ;
        RECT 42.200 24.800 42.600 25.600 ;
        RECT 43.000 24.800 43.400 25.600 ;
        RECT 45.400 25.200 45.700 26.800 ;
        RECT 45.400 24.800 45.800 25.200 ;
        RECT 46.900 25.100 47.200 26.800 ;
        RECT 47.700 26.500 48.000 27.300 ;
        RECT 47.500 26.100 48.000 26.500 ;
        RECT 47.700 25.100 48.000 26.100 ;
        RECT 39.900 23.500 40.200 24.800 ;
        RECT 40.600 23.800 41.000 24.600 ;
        RECT 44.600 23.800 45.000 24.600 ;
        RECT 45.400 23.500 45.700 24.800 ;
        RECT 46.900 24.600 47.400 25.100 ;
        RECT 47.700 24.800 49.000 25.100 ;
        RECT 39.900 23.200 41.700 23.500 ;
        RECT 39.900 23.100 40.200 23.200 ;
        RECT 36.600 21.800 38.100 22.200 ;
        RECT 37.100 21.100 38.100 21.800 ;
        RECT 39.800 21.100 40.200 23.100 ;
        RECT 41.400 23.100 41.700 23.200 ;
        RECT 43.900 23.200 45.700 23.500 ;
        RECT 43.900 23.100 44.200 23.200 ;
        RECT 41.400 21.100 41.800 23.100 ;
        RECT 43.800 21.100 44.200 23.100 ;
        RECT 45.400 23.100 45.700 23.200 ;
        RECT 45.400 21.100 45.800 23.100 ;
        RECT 47.000 21.100 47.400 24.600 ;
        RECT 48.600 21.100 49.000 24.800 ;
        RECT 51.800 21.100 52.200 29.900 ;
        RECT 54.700 28.200 55.100 29.900 ;
        RECT 54.200 27.900 55.100 28.200 ;
        RECT 55.800 27.900 56.200 29.900 ;
        RECT 56.600 28.000 57.000 29.900 ;
        RECT 58.200 28.000 58.600 29.900 ;
        RECT 59.300 28.400 59.700 29.900 ;
        RECT 56.600 27.900 58.600 28.000 ;
        RECT 59.000 27.900 59.700 28.400 ;
        RECT 61.400 27.900 61.800 29.900 ;
        RECT 53.400 26.800 53.800 27.600 ;
        RECT 54.200 26.100 54.600 27.900 ;
        RECT 55.900 27.200 56.200 27.900 ;
        RECT 56.700 27.700 58.500 27.900 ;
        RECT 57.800 27.200 58.200 27.400 ;
        RECT 55.800 26.800 57.100 27.200 ;
        RECT 57.800 26.900 58.600 27.200 ;
        RECT 58.200 26.800 58.600 26.900 ;
        RECT 56.800 26.200 57.100 26.800 ;
        RECT 54.200 25.800 56.100 26.100 ;
        RECT 56.600 25.800 57.100 26.200 ;
        RECT 57.400 26.100 57.800 26.600 ;
        RECT 59.000 26.200 59.300 27.900 ;
        RECT 61.400 27.800 61.700 27.900 ;
        RECT 62.200 27.800 62.600 28.600 ;
        RECT 60.800 27.600 61.700 27.800 ;
        RECT 59.600 27.500 61.700 27.600 ;
        RECT 59.600 27.300 61.100 27.500 ;
        RECT 59.600 27.200 60.000 27.300 ;
        RECT 58.200 26.100 58.600 26.200 ;
        RECT 57.400 25.800 58.600 26.100 ;
        RECT 59.000 25.800 59.400 26.200 ;
        RECT 54.200 21.100 54.600 25.800 ;
        RECT 55.800 25.200 56.100 25.800 ;
        RECT 55.000 24.400 55.400 25.200 ;
        RECT 55.800 25.100 56.200 25.200 ;
        RECT 56.800 25.100 57.100 25.800 ;
        RECT 59.000 25.200 59.300 25.800 ;
        RECT 59.700 25.500 60.000 27.200 ;
        RECT 61.400 27.100 61.800 27.200 ;
        RECT 63.000 27.100 63.400 29.900 ;
        RECT 64.100 28.200 64.500 29.900 ;
        RECT 64.100 27.900 65.000 28.200 ;
        RECT 66.200 27.900 66.600 29.900 ;
        RECT 67.000 28.000 67.400 29.900 ;
        RECT 68.600 28.000 69.000 29.900 ;
        RECT 70.700 29.200 71.100 29.900 ;
        RECT 73.700 29.200 74.100 29.500 ;
        RECT 70.700 28.800 71.400 29.200 ;
        RECT 73.700 28.800 74.600 29.200 ;
        RECT 70.700 28.200 71.100 28.800 ;
        RECT 67.000 27.900 69.000 28.000 ;
        RECT 70.200 27.900 71.100 28.200 ;
        RECT 73.700 28.000 74.100 28.800 ;
        RECT 75.800 28.500 76.200 29.500 ;
        RECT 61.400 26.800 63.400 27.100 ;
        RECT 61.400 26.400 61.800 26.800 ;
        RECT 59.700 25.200 60.900 25.500 ;
        RECT 55.800 24.800 56.500 25.100 ;
        RECT 56.800 24.800 57.300 25.100 ;
        RECT 56.200 24.200 56.500 24.800 ;
        RECT 56.200 23.800 56.600 24.200 ;
        RECT 56.900 21.100 57.300 24.800 ;
        RECT 59.000 21.100 59.400 25.200 ;
        RECT 60.600 23.100 60.900 25.200 ;
        RECT 60.600 21.100 61.000 23.100 ;
        RECT 63.000 21.100 63.400 26.800 ;
        RECT 63.800 24.400 64.200 25.200 ;
        RECT 64.600 21.100 65.000 27.900 ;
        RECT 65.400 26.800 65.800 27.600 ;
        RECT 66.300 27.200 66.600 27.900 ;
        RECT 67.100 27.700 68.900 27.900 ;
        RECT 68.200 27.200 68.600 27.400 ;
        RECT 66.200 26.800 67.500 27.200 ;
        RECT 68.200 26.900 69.000 27.200 ;
        RECT 68.600 26.800 69.000 26.900 ;
        RECT 69.400 26.800 69.800 27.600 ;
        RECT 66.200 26.100 66.600 26.200 ;
        RECT 67.200 26.100 67.500 26.800 ;
        RECT 66.200 25.800 67.500 26.100 ;
        RECT 67.800 25.800 68.200 26.600 ;
        RECT 65.400 25.100 65.800 25.200 ;
        RECT 66.200 25.100 66.600 25.200 ;
        RECT 67.200 25.100 67.500 25.800 ;
        RECT 65.400 24.800 66.900 25.100 ;
        RECT 67.200 24.800 67.700 25.100 ;
        RECT 66.600 24.200 66.900 24.800 ;
        RECT 66.600 23.800 67.000 24.200 ;
        RECT 67.300 21.100 67.700 24.800 ;
        RECT 70.200 21.100 70.600 27.900 ;
        RECT 73.300 27.700 74.100 28.000 ;
        RECT 73.300 27.500 73.700 27.700 ;
        RECT 73.300 27.200 73.600 27.500 ;
        RECT 75.900 27.400 76.200 28.500 ;
        RECT 72.600 26.800 73.600 27.200 ;
        RECT 74.100 27.100 76.200 27.400 ;
        RECT 77.400 28.900 77.800 29.900 ;
        RECT 77.400 27.200 77.700 28.900 ;
        RECT 78.200 27.800 78.600 28.600 ;
        RECT 79.000 27.800 79.400 28.600 ;
        RECT 74.100 26.900 74.600 27.100 ;
        RECT 71.000 26.100 71.400 26.200 ;
        RECT 72.600 26.100 73.000 26.200 ;
        RECT 71.000 25.800 73.000 26.100 ;
        RECT 72.600 25.400 73.000 25.800 ;
        RECT 71.000 24.400 71.400 25.200 ;
        RECT 73.300 24.900 73.600 26.800 ;
        RECT 73.900 26.500 74.600 26.900 ;
        RECT 77.400 26.800 77.800 27.200 ;
        RECT 74.300 25.500 74.600 26.500 ;
        RECT 75.000 25.800 75.400 26.600 ;
        RECT 75.800 25.800 76.200 26.600 ;
        RECT 74.300 25.200 76.200 25.500 ;
        RECT 76.600 25.400 77.000 26.200 ;
        RECT 73.300 24.600 74.100 24.900 ;
        RECT 73.700 21.100 74.100 24.600 ;
        RECT 75.900 23.500 76.200 25.200 ;
        RECT 77.400 25.100 77.700 26.800 ;
        RECT 75.800 21.500 76.200 23.500 ;
        RECT 76.900 24.700 77.800 25.100 ;
        RECT 76.900 22.200 77.300 24.700 ;
        RECT 76.900 21.800 77.800 22.200 ;
        RECT 76.900 21.100 77.300 21.800 ;
        RECT 79.800 21.100 80.200 29.900 ;
        RECT 82.200 27.900 82.600 29.900 ;
        RECT 82.900 28.200 83.300 28.600 ;
        RECT 81.400 26.400 81.800 27.200 ;
        RECT 80.600 26.100 81.000 26.200 ;
        RECT 82.200 26.100 82.500 27.900 ;
        RECT 83.000 27.800 83.400 28.200 ;
        RECT 83.800 28.000 84.200 29.900 ;
        RECT 85.400 28.000 85.800 29.900 ;
        RECT 83.800 27.900 85.800 28.000 ;
        RECT 86.200 27.900 86.600 29.900 ;
        RECT 87.000 27.900 87.400 29.900 ;
        RECT 87.800 28.000 88.200 29.900 ;
        RECT 89.400 28.000 89.800 29.900 ;
        RECT 87.800 27.900 89.800 28.000 ;
        RECT 83.900 27.700 85.700 27.900 ;
        RECT 84.200 27.200 84.600 27.400 ;
        RECT 86.200 27.200 86.500 27.900 ;
        RECT 87.100 27.200 87.400 27.900 ;
        RECT 87.900 27.700 89.700 27.900 ;
        RECT 89.000 27.200 89.400 27.400 ;
        RECT 83.800 26.900 84.600 27.200 ;
        RECT 83.800 26.800 84.200 26.900 ;
        RECT 85.300 26.800 86.600 27.200 ;
        RECT 87.000 26.800 88.300 27.200 ;
        RECT 89.000 27.100 89.800 27.200 ;
        RECT 90.200 27.100 90.600 29.900 ;
        RECT 92.600 28.900 93.000 29.900 ;
        RECT 91.000 28.100 91.400 28.600 ;
        RECT 92.600 28.100 92.900 28.900 ;
        RECT 91.000 27.800 92.900 28.100 ;
        RECT 93.400 27.800 93.800 28.600 ;
        RECT 95.800 27.900 96.200 29.900 ;
        RECT 96.500 28.200 96.900 28.600 ;
        RECT 98.700 28.200 99.100 29.900 ;
        RECT 89.000 26.900 90.600 27.100 ;
        RECT 89.400 26.800 90.600 26.900 ;
        RECT 83.000 26.100 83.400 26.200 ;
        RECT 80.600 25.800 81.400 26.100 ;
        RECT 82.200 25.800 83.400 26.100 ;
        RECT 81.000 25.600 81.400 25.800 ;
        RECT 83.000 25.100 83.300 25.800 ;
        RECT 85.300 25.100 85.600 26.800 ;
        RECT 86.200 25.100 86.600 25.200 ;
        RECT 80.600 24.800 82.600 25.100 ;
        RECT 80.600 21.100 81.000 24.800 ;
        RECT 82.200 21.100 82.600 24.800 ;
        RECT 83.000 21.100 83.400 25.100 ;
        RECT 85.100 24.800 85.600 25.100 ;
        RECT 85.900 24.800 86.600 25.100 ;
        RECT 87.000 25.100 87.400 25.200 ;
        RECT 88.000 25.100 88.300 26.800 ;
        RECT 88.600 26.100 89.000 26.600 ;
        RECT 89.400 26.100 89.800 26.200 ;
        RECT 88.600 25.800 89.800 26.100 ;
        RECT 87.000 24.800 87.700 25.100 ;
        RECT 88.000 24.800 88.500 25.100 ;
        RECT 85.100 21.100 85.500 24.800 ;
        RECT 85.900 24.200 86.200 24.800 ;
        RECT 85.800 23.800 86.200 24.200 ;
        RECT 87.400 24.200 87.700 24.800 ;
        RECT 87.400 23.800 87.800 24.200 ;
        RECT 88.100 21.100 88.500 24.800 ;
        RECT 90.200 21.100 90.600 26.800 ;
        RECT 92.600 27.200 92.900 27.800 ;
        RECT 92.600 26.800 93.000 27.200 ;
        RECT 92.600 26.200 92.900 26.800 ;
        RECT 95.000 26.400 95.400 27.200 ;
        RECT 91.800 25.400 92.200 26.200 ;
        RECT 92.600 25.800 93.000 26.200 ;
        RECT 94.200 26.100 94.600 26.200 ;
        RECT 95.800 26.100 96.100 27.900 ;
        RECT 96.600 27.800 97.000 28.200 ;
        RECT 98.200 27.900 99.100 28.200 ;
        RECT 101.400 27.900 101.800 29.900 ;
        RECT 103.500 29.200 103.900 29.900 ;
        RECT 103.500 28.800 104.200 29.200 ;
        RECT 103.500 28.400 103.900 28.800 ;
        RECT 103.500 27.900 104.200 28.400 ;
        RECT 97.400 26.800 97.800 27.600 ;
        RECT 98.200 27.100 98.600 27.900 ;
        RECT 101.500 27.800 101.800 27.900 ;
        RECT 101.500 27.600 102.400 27.800 ;
        RECT 101.500 27.500 103.600 27.600 ;
        RECT 102.100 27.300 103.600 27.500 ;
        RECT 103.200 27.200 103.600 27.300 ;
        RECT 99.800 27.100 100.200 27.200 ;
        RECT 98.200 26.800 100.200 27.100 ;
        RECT 96.600 26.100 97.000 26.200 ;
        RECT 94.200 25.800 95.000 26.100 ;
        RECT 95.800 25.800 97.000 26.100 ;
        RECT 92.600 25.100 92.900 25.800 ;
        RECT 94.600 25.600 95.000 25.800 ;
        RECT 96.600 25.100 96.900 25.800 ;
        RECT 92.100 24.700 93.000 25.100 ;
        RECT 94.200 24.800 96.200 25.100 ;
        RECT 92.100 21.100 92.500 24.700 ;
        RECT 94.200 21.100 94.600 24.800 ;
        RECT 95.800 21.100 96.200 24.800 ;
        RECT 96.600 21.100 97.000 25.100 ;
        RECT 98.200 21.100 98.600 26.800 ;
        RECT 101.400 26.400 101.800 27.200 ;
        RECT 102.200 26.600 102.800 27.000 ;
        RECT 102.300 26.200 102.600 26.600 ;
        RECT 102.200 25.800 102.600 26.200 ;
        RECT 103.200 25.500 103.500 27.200 ;
        RECT 103.900 26.200 104.200 27.900 ;
        RECT 103.800 25.800 104.200 26.200 ;
        RECT 102.300 25.200 103.500 25.500 ;
        RECT 99.000 24.400 99.400 25.200 ;
        RECT 102.300 23.100 102.600 25.200 ;
        RECT 103.900 25.100 104.200 25.800 ;
        RECT 102.200 21.100 102.600 23.100 ;
        RECT 103.800 21.100 104.200 25.100 ;
        RECT 104.600 21.100 105.000 29.900 ;
        RECT 105.400 27.800 105.800 28.600 ;
        RECT 106.200 27.900 106.600 29.900 ;
        RECT 107.000 28.000 107.400 29.900 ;
        RECT 108.600 28.000 109.000 29.900 ;
        RECT 107.000 27.900 109.000 28.000 ;
        RECT 111.000 27.900 111.400 29.900 ;
        RECT 111.700 28.200 112.100 28.600 ;
        RECT 106.300 27.200 106.600 27.900 ;
        RECT 107.100 27.700 108.900 27.900 ;
        RECT 108.200 27.200 108.600 27.400 ;
        RECT 106.200 26.800 107.500 27.200 ;
        RECT 108.200 26.900 109.000 27.200 ;
        RECT 108.600 26.800 109.000 26.900 ;
        RECT 107.200 25.200 107.500 26.800 ;
        RECT 107.800 25.800 108.200 26.600 ;
        RECT 110.200 26.400 110.600 27.200 ;
        RECT 109.400 26.100 109.800 26.200 ;
        RECT 111.000 26.100 111.300 27.900 ;
        RECT 111.800 27.800 112.200 28.200 ;
        RECT 114.200 27.800 114.600 29.900 ;
        RECT 114.900 28.200 115.300 28.600 ;
        RECT 115.000 27.800 115.400 28.200 ;
        RECT 117.400 27.900 117.800 29.900 ;
        RECT 118.100 28.200 118.500 28.600 ;
        RECT 113.400 26.400 113.800 27.200 ;
        RECT 111.800 26.100 112.200 26.200 ;
        RECT 109.400 25.800 110.200 26.100 ;
        RECT 111.000 25.800 112.200 26.100 ;
        RECT 112.600 26.100 113.000 26.200 ;
        RECT 114.200 26.100 114.500 27.800 ;
        RECT 116.600 26.400 117.000 27.200 ;
        RECT 115.000 26.100 115.400 26.200 ;
        RECT 112.600 25.800 113.400 26.100 ;
        RECT 114.200 25.800 115.400 26.100 ;
        RECT 115.800 26.100 116.200 26.200 ;
        RECT 117.400 26.100 117.700 27.900 ;
        RECT 118.200 27.800 118.600 28.200 ;
        RECT 119.000 27.900 119.400 29.900 ;
        RECT 119.800 28.000 120.200 29.900 ;
        RECT 121.400 28.000 121.800 29.900 ;
        RECT 119.800 27.900 121.800 28.000 ;
        RECT 122.200 27.900 122.600 29.900 ;
        RECT 123.000 28.000 123.400 29.900 ;
        RECT 124.600 28.000 125.000 29.900 ;
        RECT 123.000 27.900 125.000 28.000 ;
        RECT 125.400 27.900 125.800 29.900 ;
        RECT 127.500 28.400 127.900 29.900 ;
        RECT 127.500 27.900 128.200 28.400 ;
        RECT 129.900 28.200 130.300 29.900 ;
        RECT 119.100 27.200 119.400 27.900 ;
        RECT 119.900 27.700 121.700 27.900 ;
        RECT 121.000 27.200 121.400 27.400 ;
        RECT 122.300 27.200 122.600 27.900 ;
        RECT 123.100 27.700 124.900 27.900 ;
        RECT 125.500 27.800 125.800 27.900 ;
        RECT 125.500 27.600 126.400 27.800 ;
        RECT 125.500 27.500 127.600 27.600 ;
        RECT 124.200 27.200 124.600 27.400 ;
        RECT 126.100 27.300 127.600 27.500 ;
        RECT 127.200 27.200 127.600 27.300 ;
        RECT 118.200 27.100 118.600 27.200 ;
        RECT 119.000 27.100 120.300 27.200 ;
        RECT 118.200 26.800 120.300 27.100 ;
        RECT 121.000 26.900 121.800 27.200 ;
        RECT 121.400 26.800 121.800 26.900 ;
        RECT 122.200 26.800 123.500 27.200 ;
        RECT 124.200 27.100 125.000 27.200 ;
        RECT 125.400 27.100 125.800 27.200 ;
        RECT 124.200 26.900 125.800 27.100 ;
        RECT 126.400 26.900 126.800 27.000 ;
        RECT 124.600 26.800 125.800 26.900 ;
        RECT 118.200 26.100 118.600 26.200 ;
        RECT 115.800 25.800 116.600 26.100 ;
        RECT 117.400 25.800 118.600 26.100 ;
        RECT 109.800 25.600 110.200 25.800 ;
        RECT 105.400 25.100 105.800 25.200 ;
        RECT 106.200 25.100 106.600 25.200 ;
        RECT 105.400 24.800 106.900 25.100 ;
        RECT 107.200 24.800 108.200 25.200 ;
        RECT 111.800 25.100 112.100 25.800 ;
        RECT 113.000 25.600 113.400 25.800 ;
        RECT 115.000 25.100 115.300 25.800 ;
        RECT 116.200 25.600 116.600 25.800 ;
        RECT 118.200 25.100 118.500 25.800 ;
        RECT 119.000 25.100 119.400 25.200 ;
        RECT 120.000 25.100 120.300 26.800 ;
        RECT 120.600 26.100 121.000 26.600 ;
        RECT 123.200 26.100 123.500 26.800 ;
        RECT 120.600 25.800 123.500 26.100 ;
        RECT 123.800 25.800 124.200 26.600 ;
        RECT 125.400 26.400 125.800 26.800 ;
        RECT 126.300 26.600 126.800 26.900 ;
        RECT 126.300 26.200 126.600 26.600 ;
        RECT 126.200 25.800 126.600 26.200 ;
        RECT 122.200 25.100 122.600 25.200 ;
        RECT 123.200 25.100 123.500 25.800 ;
        RECT 127.200 25.500 127.500 27.200 ;
        RECT 127.900 26.200 128.200 27.900 ;
        RECT 129.400 27.900 130.300 28.200 ;
        RECT 131.800 28.900 132.200 29.900 ;
        RECT 128.600 26.800 129.000 27.600 ;
        RECT 129.400 27.100 129.800 27.900 ;
        RECT 131.800 27.200 132.100 28.900 ;
        RECT 132.600 27.800 133.000 28.600 ;
        RECT 133.400 28.000 133.800 29.900 ;
        RECT 135.000 28.000 135.400 29.900 ;
        RECT 133.400 27.900 135.400 28.000 ;
        RECT 135.800 27.900 136.200 29.900 ;
        RECT 138.200 27.900 138.600 29.900 ;
        RECT 138.900 28.200 139.300 28.600 ;
        RECT 133.500 27.700 135.300 27.900 ;
        RECT 133.800 27.200 134.200 27.400 ;
        RECT 135.800 27.200 136.100 27.900 ;
        RECT 130.200 27.100 130.600 27.200 ;
        RECT 129.400 26.800 130.600 27.100 ;
        RECT 131.800 26.800 132.200 27.200 ;
        RECT 133.400 26.900 134.200 27.200 ;
        RECT 133.400 26.800 133.800 26.900 ;
        RECT 134.900 26.800 136.200 27.200 ;
        RECT 127.800 25.800 128.200 26.200 ;
        RECT 126.300 25.200 127.500 25.500 ;
        RECT 109.400 24.800 111.400 25.100 ;
        RECT 106.600 24.200 106.900 24.800 ;
        RECT 106.600 23.800 107.000 24.200 ;
        RECT 107.300 21.100 107.700 24.800 ;
        RECT 109.400 21.100 109.800 24.800 ;
        RECT 111.000 21.100 111.400 24.800 ;
        RECT 111.800 21.100 112.200 25.100 ;
        RECT 112.600 24.800 114.600 25.100 ;
        RECT 112.600 21.100 113.000 24.800 ;
        RECT 114.200 21.100 114.600 24.800 ;
        RECT 115.000 21.100 115.400 25.100 ;
        RECT 115.800 24.800 117.800 25.100 ;
        RECT 115.800 21.100 116.200 24.800 ;
        RECT 117.400 21.100 117.800 24.800 ;
        RECT 118.200 21.100 118.600 25.100 ;
        RECT 119.000 24.800 119.700 25.100 ;
        RECT 120.000 24.800 120.500 25.100 ;
        RECT 122.200 24.800 122.900 25.100 ;
        RECT 123.200 24.800 123.700 25.100 ;
        RECT 119.400 24.200 119.700 24.800 ;
        RECT 119.400 23.800 119.800 24.200 ;
        RECT 120.100 21.100 120.500 24.800 ;
        RECT 122.600 24.200 122.900 24.800 ;
        RECT 122.600 23.800 123.000 24.200 ;
        RECT 123.300 21.100 123.700 24.800 ;
        RECT 126.300 23.100 126.600 25.200 ;
        RECT 127.900 25.100 128.200 25.800 ;
        RECT 126.200 21.100 126.600 23.100 ;
        RECT 127.800 21.100 128.200 25.100 ;
        RECT 129.400 21.100 129.800 26.800 ;
        RECT 131.000 25.400 131.400 26.200 ;
        RECT 130.200 24.100 130.600 25.200 ;
        RECT 131.800 25.100 132.100 26.800 ;
        RECT 132.600 26.100 133.000 26.200 ;
        RECT 134.200 26.100 134.600 26.600 ;
        RECT 132.600 25.800 134.600 26.100 ;
        RECT 134.900 26.100 135.200 26.800 ;
        RECT 137.400 26.400 137.800 27.200 ;
        RECT 136.600 26.100 137.000 26.200 ;
        RECT 138.200 26.100 138.500 27.900 ;
        RECT 139.000 27.800 139.400 28.200 ;
        RECT 139.000 26.100 139.400 26.200 ;
        RECT 134.900 25.800 137.400 26.100 ;
        RECT 138.200 25.800 139.400 26.100 ;
        RECT 134.900 25.100 135.200 25.800 ;
        RECT 137.000 25.600 137.400 25.800 ;
        RECT 135.800 25.100 136.200 25.200 ;
        RECT 139.000 25.100 139.300 25.800 ;
        RECT 131.300 24.700 132.200 25.100 ;
        RECT 134.700 24.800 135.200 25.100 ;
        RECT 135.500 24.800 136.200 25.100 ;
        RECT 136.600 24.800 138.600 25.100 ;
        RECT 131.300 24.100 131.700 24.700 ;
        RECT 130.200 23.800 131.700 24.100 ;
        RECT 131.300 21.100 131.700 23.800 ;
        RECT 134.700 21.100 135.100 24.800 ;
        RECT 135.500 24.200 135.800 24.800 ;
        RECT 135.400 23.800 135.800 24.200 ;
        RECT 136.600 21.100 137.000 24.800 ;
        RECT 138.200 21.100 138.600 24.800 ;
        RECT 139.000 21.100 139.400 25.100 ;
        RECT 140.600 21.100 141.000 29.900 ;
        RECT 141.400 26.800 141.800 27.600 ;
        RECT 141.400 26.100 141.800 26.200 ;
        RECT 142.200 26.100 142.600 29.900 ;
        RECT 144.600 28.900 145.000 29.900 ;
        RECT 143.000 27.100 143.400 27.600 ;
        RECT 144.700 27.200 145.000 28.900 ;
        RECT 147.000 28.900 147.400 29.900 ;
        RECT 149.400 29.100 149.800 29.900 ;
        RECT 150.200 29.100 150.600 29.200 ;
        RECT 144.600 27.100 145.000 27.200 ;
        RECT 143.000 26.800 145.000 27.100 ;
        RECT 145.400 27.800 145.800 28.200 ;
        RECT 145.400 27.100 145.700 27.800 ;
        RECT 147.000 27.200 147.300 28.900 ;
        RECT 149.400 28.800 150.600 29.100 ;
        RECT 147.800 27.800 148.200 28.600 ;
        RECT 147.000 27.100 147.400 27.200 ;
        RECT 145.400 26.800 147.400 27.100 ;
        RECT 141.400 25.800 142.600 26.100 ;
        RECT 142.200 21.100 142.600 25.800 ;
        RECT 144.700 25.100 145.000 26.800 ;
        RECT 145.400 26.100 145.800 26.200 ;
        RECT 146.200 26.100 146.600 26.200 ;
        RECT 145.400 25.800 146.600 26.100 ;
        RECT 145.400 25.400 145.800 25.800 ;
        RECT 146.200 25.400 146.600 25.800 ;
        RECT 147.000 25.100 147.300 26.800 ;
        RECT 144.600 24.700 145.500 25.100 ;
        RECT 145.100 21.100 145.500 24.700 ;
        RECT 146.500 24.700 147.400 25.100 ;
        RECT 146.500 21.100 146.900 24.700 ;
        RECT 149.400 21.100 149.800 28.800 ;
        RECT 0.600 17.900 1.000 19.900 ;
        RECT 0.700 17.800 1.000 17.900 ;
        RECT 2.200 17.900 2.600 19.900 ;
        RECT 3.800 17.900 4.200 19.900 ;
        RECT 2.200 17.800 2.500 17.900 ;
        RECT 0.700 17.500 2.500 17.800 ;
        RECT 3.900 17.800 4.200 17.900 ;
        RECT 5.400 17.900 5.800 19.900 ;
        RECT 8.100 19.200 8.500 19.900 ;
        RECT 8.100 18.800 9.000 19.200 ;
        RECT 5.400 17.800 5.700 17.900 ;
        RECT 3.900 17.500 5.700 17.800 ;
        RECT 0.700 16.200 1.000 17.500 ;
        RECT 1.400 16.400 1.800 17.200 ;
        RECT 3.900 16.200 4.200 17.500 ;
        RECT 4.600 16.400 5.000 17.200 ;
        RECT 7.400 16.800 7.800 17.200 ;
        RECT 7.400 16.200 7.700 16.800 ;
        RECT 8.100 16.200 8.500 18.800 ;
        RECT 0.600 15.800 1.000 16.200 ;
        RECT 0.700 14.200 1.000 15.800 ;
        RECT 3.000 15.400 3.400 16.200 ;
        RECT 3.800 15.800 4.200 16.200 ;
        RECT 3.900 15.200 4.200 15.800 ;
        RECT 6.200 15.400 6.600 16.200 ;
        RECT 7.000 15.900 7.700 16.200 ;
        RECT 8.000 15.900 8.500 16.200 ;
        RECT 10.200 15.900 10.600 19.900 ;
        RECT 11.000 16.200 11.400 19.900 ;
        RECT 12.600 16.200 13.000 19.900 ;
        RECT 14.500 18.200 14.900 19.900 ;
        RECT 14.500 17.800 15.400 18.200 ;
        RECT 13.800 16.800 14.200 17.200 ;
        RECT 13.800 16.200 14.100 16.800 ;
        RECT 14.500 16.200 14.900 17.800 ;
        RECT 11.000 15.900 13.000 16.200 ;
        RECT 13.400 15.900 14.100 16.200 ;
        RECT 14.400 15.900 14.900 16.200 ;
        RECT 17.900 16.200 18.300 19.900 ;
        RECT 19.800 17.900 20.200 19.900 ;
        RECT 19.900 17.800 20.200 17.900 ;
        RECT 21.400 17.900 21.800 19.900 ;
        RECT 21.400 17.800 21.700 17.900 ;
        RECT 19.900 17.500 21.700 17.800 ;
        RECT 23.800 17.800 24.200 19.900 ;
        RECT 25.400 17.900 25.800 19.900 ;
        RECT 25.400 17.800 25.700 17.900 ;
        RECT 23.800 17.500 25.700 17.800 ;
        RECT 18.600 16.800 19.000 17.200 ;
        RECT 18.700 16.200 19.000 16.800 ;
        RECT 19.900 16.200 20.200 17.500 ;
        RECT 20.600 16.400 21.000 17.200 ;
        RECT 23.800 17.100 24.100 17.500 ;
        RECT 22.200 16.800 24.100 17.100 ;
        RECT 17.900 15.900 18.400 16.200 ;
        RECT 18.700 15.900 19.400 16.200 ;
        RECT 7.000 15.800 7.400 15.900 ;
        RECT 1.800 14.800 2.600 15.200 ;
        RECT 3.800 14.800 4.200 15.200 ;
        RECT 5.000 14.800 5.800 15.200 ;
        RECT 3.900 14.200 4.200 14.800 ;
        RECT 8.000 14.200 8.300 15.900 ;
        RECT 10.300 15.200 10.600 15.900 ;
        RECT 13.400 15.800 13.800 15.900 ;
        RECT 12.200 15.200 12.600 15.400 ;
        RECT 8.600 15.100 9.000 15.200 ;
        RECT 10.200 15.100 11.400 15.200 ;
        RECT 8.600 14.900 11.400 15.100 ;
        RECT 12.200 14.900 13.000 15.200 ;
        RECT 8.600 14.800 10.600 14.900 ;
        RECT 8.600 14.400 9.000 14.800 ;
        RECT 0.700 14.100 1.500 14.200 ;
        RECT 3.900 14.100 4.700 14.200 ;
        RECT 0.700 13.900 1.600 14.100 ;
        RECT 3.900 13.900 4.800 14.100 ;
        RECT 1.200 11.100 1.600 13.900 ;
        RECT 4.400 11.100 4.800 13.900 ;
        RECT 7.000 13.800 8.300 14.200 ;
        RECT 9.400 14.100 9.800 14.200 ;
        RECT 9.000 13.800 9.800 14.100 ;
        RECT 7.100 13.100 7.400 13.800 ;
        RECT 9.000 13.600 9.400 13.800 ;
        RECT 7.900 13.100 9.700 13.300 ;
        RECT 7.000 11.100 7.400 13.100 ;
        RECT 7.800 13.000 9.800 13.100 ;
        RECT 7.800 11.100 8.200 13.000 ;
        RECT 9.400 11.100 9.800 13.000 ;
        RECT 10.200 12.800 10.600 13.200 ;
        RECT 11.100 13.100 11.400 14.900 ;
        RECT 12.600 14.800 13.000 14.900 ;
        RECT 11.800 13.800 12.200 14.600 ;
        RECT 14.400 14.200 14.700 15.900 ;
        RECT 18.100 15.200 18.400 15.900 ;
        RECT 19.000 15.800 19.400 15.900 ;
        RECT 19.800 15.800 20.200 16.200 ;
        RECT 15.000 15.100 15.400 15.200 ;
        RECT 17.400 15.100 17.800 15.200 ;
        RECT 15.000 14.800 17.800 15.100 ;
        RECT 15.000 14.400 15.400 14.800 ;
        RECT 17.400 14.400 17.800 14.800 ;
        RECT 18.100 14.800 18.600 15.200 ;
        RECT 18.100 14.200 18.400 14.800 ;
        RECT 19.900 14.200 20.200 15.800 ;
        RECT 22.200 16.200 22.500 16.800 ;
        RECT 24.600 16.400 25.000 17.200 ;
        RECT 25.400 16.200 25.700 17.500 ;
        RECT 22.200 15.400 22.600 16.200 ;
        RECT 23.000 15.400 23.400 16.200 ;
        RECT 25.400 15.800 25.800 16.200 ;
        RECT 26.200 15.900 26.600 19.900 ;
        RECT 27.000 16.200 27.400 19.900 ;
        RECT 28.600 16.200 29.000 19.900 ;
        RECT 27.000 15.900 29.000 16.200 ;
        RECT 21.000 14.800 21.800 15.200 ;
        RECT 23.800 14.800 24.600 15.200 ;
        RECT 25.400 14.200 25.700 15.800 ;
        RECT 26.300 15.200 26.600 15.900 ;
        RECT 28.200 15.200 28.600 15.400 ;
        RECT 26.200 14.900 27.400 15.200 ;
        RECT 28.200 14.900 29.000 15.200 ;
        RECT 26.200 14.800 26.600 14.900 ;
        RECT 13.400 13.800 14.700 14.200 ;
        RECT 15.800 14.100 16.200 14.200 ;
        RECT 16.600 14.100 17.000 14.200 ;
        RECT 15.400 13.800 17.400 14.100 ;
        RECT 18.100 13.800 19.400 14.200 ;
        RECT 19.900 14.100 20.700 14.200 ;
        RECT 24.900 14.100 25.700 14.200 ;
        RECT 19.900 13.900 20.800 14.100 ;
        RECT 13.500 13.100 13.800 13.800 ;
        RECT 15.400 13.600 15.800 13.800 ;
        RECT 17.000 13.600 17.400 13.800 ;
        RECT 14.300 13.100 16.100 13.300 ;
        RECT 16.700 13.100 18.500 13.300 ;
        RECT 19.000 13.100 19.300 13.800 ;
        RECT 10.300 12.400 10.700 12.800 ;
        RECT 11.000 11.100 11.400 13.100 ;
        RECT 13.400 11.100 13.800 13.100 ;
        RECT 14.200 13.000 16.200 13.100 ;
        RECT 14.200 11.100 14.600 13.000 ;
        RECT 15.800 11.100 16.200 13.000 ;
        RECT 16.600 13.000 18.600 13.100 ;
        RECT 16.600 11.100 17.000 13.000 ;
        RECT 18.200 11.100 18.600 13.000 ;
        RECT 19.000 11.100 19.400 13.100 ;
        RECT 20.400 11.100 20.800 13.900 ;
        RECT 24.800 13.900 25.700 14.100 ;
        RECT 24.800 11.100 25.200 13.900 ;
        RECT 26.200 12.800 26.600 13.200 ;
        RECT 27.100 13.100 27.400 14.900 ;
        RECT 28.600 14.800 29.000 14.900 ;
        RECT 27.800 13.800 28.200 14.600 ;
        RECT 29.400 13.400 29.800 14.200 ;
        RECT 26.300 12.400 26.700 12.800 ;
        RECT 27.000 11.100 27.400 13.100 ;
        RECT 30.200 13.100 30.600 19.900 ;
        RECT 32.600 17.900 33.000 19.900 ;
        RECT 31.000 15.800 31.400 16.600 ;
        RECT 32.700 15.800 33.000 17.900 ;
        RECT 34.200 15.900 34.600 19.900 ;
        RECT 35.000 17.900 35.400 19.900 ;
        RECT 35.100 17.800 35.400 17.900 ;
        RECT 36.600 17.900 37.000 19.900 ;
        RECT 36.600 17.800 36.900 17.900 ;
        RECT 35.100 17.500 36.900 17.800 ;
        RECT 35.100 16.200 35.400 17.500 ;
        RECT 35.800 16.400 36.200 17.200 ;
        RECT 32.700 15.500 33.900 15.800 ;
        RECT 32.600 14.800 33.000 15.200 ;
        RECT 31.800 13.800 32.200 14.600 ;
        RECT 32.700 14.400 33.000 14.800 ;
        RECT 32.700 14.100 33.200 14.400 ;
        RECT 32.800 14.000 33.200 14.100 ;
        RECT 33.600 13.800 33.900 15.500 ;
        RECT 34.300 15.200 34.600 15.900 ;
        RECT 35.000 15.800 35.400 16.200 ;
        RECT 35.100 15.200 35.400 15.800 ;
        RECT 37.400 15.400 37.800 16.200 ;
        RECT 38.200 15.900 38.600 19.900 ;
        RECT 39.000 16.200 39.400 19.900 ;
        RECT 40.600 16.200 41.000 19.900 ;
        RECT 39.000 15.900 41.000 16.200 ;
        RECT 38.300 15.200 38.600 15.900 ;
        RECT 40.200 15.200 40.600 15.400 ;
        RECT 34.200 14.800 34.600 15.200 ;
        RECT 35.000 14.800 35.400 15.200 ;
        RECT 36.200 14.800 37.000 15.200 ;
        RECT 38.200 14.900 39.400 15.200 ;
        RECT 40.200 14.900 41.000 15.200 ;
        RECT 38.200 14.800 38.600 14.900 ;
        RECT 33.600 13.700 34.000 13.800 ;
        RECT 32.500 13.500 34.000 13.700 ;
        RECT 31.900 13.400 34.000 13.500 ;
        RECT 31.900 13.200 32.800 13.400 ;
        RECT 31.900 13.100 32.200 13.200 ;
        RECT 34.300 13.100 34.600 14.800 ;
        RECT 35.100 14.200 35.400 14.800 ;
        RECT 35.100 14.100 35.900 14.200 ;
        RECT 35.100 13.900 36.000 14.100 ;
        RECT 30.200 12.800 31.100 13.100 ;
        RECT 30.700 12.200 31.100 12.800 ;
        RECT 30.200 11.800 31.100 12.200 ;
        RECT 30.700 11.100 31.100 11.800 ;
        RECT 31.800 11.100 32.200 13.100 ;
        RECT 33.900 12.600 34.600 13.100 ;
        RECT 33.900 11.100 34.300 12.600 ;
        RECT 35.600 11.100 36.000 13.900 ;
        RECT 38.200 12.800 38.600 13.200 ;
        RECT 39.100 13.100 39.400 14.900 ;
        RECT 40.600 14.800 41.000 14.900 ;
        RECT 39.800 13.800 40.200 14.600 ;
        RECT 41.400 14.100 41.800 14.200 ;
        RECT 42.200 14.100 42.600 19.900 ;
        RECT 43.000 16.200 43.400 19.900 ;
        RECT 44.600 16.400 45.000 19.900 ;
        RECT 43.000 15.900 44.300 16.200 ;
        RECT 44.600 15.900 45.100 16.400 ;
        RECT 46.200 15.900 46.600 19.900 ;
        RECT 47.000 16.200 47.400 19.900 ;
        RECT 48.600 16.200 49.000 19.900 ;
        RECT 47.000 15.900 49.000 16.200 ;
        RECT 51.000 16.200 51.400 19.900 ;
        RECT 52.600 16.200 53.000 19.900 ;
        RECT 51.000 15.900 53.000 16.200 ;
        RECT 53.400 15.900 53.800 19.900 ;
        RECT 54.200 16.200 54.600 19.900 ;
        RECT 55.800 16.400 56.200 19.900 ;
        RECT 59.300 19.200 59.700 19.900 ;
        RECT 59.300 18.800 60.200 19.200 ;
        RECT 59.300 16.400 59.700 18.800 ;
        RECT 61.400 17.500 61.800 19.500 ;
        RECT 54.200 15.900 55.500 16.200 ;
        RECT 41.400 13.800 42.600 14.100 ;
        RECT 38.300 12.400 38.700 12.800 ;
        RECT 39.000 11.100 39.400 13.100 ;
        RECT 41.400 12.400 41.800 13.200 ;
        RECT 42.200 11.100 42.600 13.800 ;
        RECT 44.000 14.900 44.300 15.900 ;
        RECT 44.000 14.500 44.500 14.900 ;
        RECT 44.000 13.700 44.300 14.500 ;
        RECT 44.800 14.200 45.100 15.900 ;
        RECT 46.300 15.200 46.600 15.900 ;
        RECT 48.200 15.200 48.600 15.400 ;
        RECT 51.400 15.200 51.800 15.400 ;
        RECT 53.400 15.200 53.700 15.900 ;
        RECT 46.200 14.900 47.400 15.200 ;
        RECT 48.200 14.900 49.000 15.200 ;
        RECT 46.200 14.800 46.600 14.900 ;
        RECT 44.600 14.100 45.100 14.200 ;
        RECT 45.400 14.100 45.800 14.200 ;
        RECT 44.600 13.800 45.800 14.100 ;
        RECT 43.000 13.400 44.300 13.700 ;
        RECT 43.000 11.100 43.400 13.400 ;
        RECT 44.800 13.100 45.100 13.800 ;
        RECT 44.600 12.800 45.100 13.100 ;
        RECT 46.200 12.800 46.600 13.200 ;
        RECT 47.100 13.100 47.400 14.900 ;
        RECT 48.600 14.800 49.000 14.900 ;
        RECT 51.000 14.900 51.800 15.200 ;
        RECT 52.600 14.900 53.800 15.200 ;
        RECT 51.000 14.800 51.400 14.900 ;
        RECT 44.600 11.100 45.000 12.800 ;
        RECT 46.300 12.400 46.700 12.800 ;
        RECT 47.000 11.100 47.400 13.100 ;
        RECT 52.600 13.100 52.900 14.900 ;
        RECT 53.400 14.800 53.800 14.900 ;
        RECT 55.200 14.900 55.500 15.900 ;
        RECT 55.800 15.800 56.300 16.400 ;
        RECT 55.200 14.500 55.700 14.900 ;
        RECT 55.200 13.700 55.500 14.500 ;
        RECT 56.000 14.200 56.300 15.800 ;
        RECT 58.900 16.100 59.700 16.400 ;
        RECT 58.900 14.200 59.200 16.100 ;
        RECT 61.500 15.800 61.800 17.500 ;
        RECT 59.900 15.500 61.800 15.800 ;
        RECT 59.900 14.500 60.200 15.500 ;
        RECT 55.800 13.800 56.300 14.200 ;
        RECT 58.200 13.800 59.200 14.200 ;
        RECT 59.500 14.100 60.200 14.500 ;
        RECT 61.400 14.400 61.800 15.200 ;
        RECT 63.000 15.100 63.400 19.900 ;
        RECT 64.100 16.300 64.500 19.900 ;
        RECT 64.100 15.900 65.000 16.300 ;
        RECT 63.800 15.100 64.200 15.600 ;
        RECT 63.000 14.800 64.200 15.100 ;
        RECT 54.200 13.400 55.500 13.700 ;
        RECT 52.600 11.100 53.000 13.100 ;
        RECT 53.400 12.800 53.800 13.200 ;
        RECT 53.300 12.400 53.700 12.800 ;
        RECT 54.200 11.100 54.600 13.400 ;
        RECT 56.000 13.100 56.300 13.800 ;
        RECT 55.800 12.800 56.300 13.100 ;
        RECT 58.900 13.500 59.200 13.800 ;
        RECT 59.700 13.900 60.200 14.100 ;
        RECT 59.700 13.600 61.800 13.900 ;
        RECT 58.900 13.300 59.300 13.500 ;
        RECT 58.900 13.000 59.700 13.300 ;
        RECT 55.800 11.100 56.200 12.800 ;
        RECT 59.300 11.500 59.700 13.000 ;
        RECT 61.500 12.500 61.800 13.600 ;
        RECT 61.400 11.500 61.800 12.500 ;
        RECT 63.000 11.100 63.400 14.800 ;
        RECT 64.600 14.200 64.900 15.900 ;
        RECT 64.600 13.800 65.000 14.200 ;
        RECT 63.800 13.100 64.200 13.200 ;
        RECT 64.600 13.100 64.900 13.800 ;
        RECT 63.800 12.800 64.900 13.100 ;
        RECT 64.600 12.100 64.900 12.800 ;
        RECT 65.400 12.400 65.800 13.200 ;
        RECT 64.600 11.100 65.000 12.100 ;
        RECT 67.000 11.100 67.400 19.900 ;
        RECT 68.100 16.300 68.500 19.900 ;
        RECT 68.100 15.900 69.000 16.300 ;
        RECT 71.500 16.200 71.900 19.900 ;
        RECT 74.200 17.800 74.600 19.900 ;
        RECT 75.800 17.900 76.200 19.900 ;
        RECT 75.800 17.800 76.100 17.900 ;
        RECT 74.300 17.500 76.100 17.800 ;
        RECT 72.200 16.800 72.600 17.200 ;
        RECT 74.200 17.100 74.600 17.200 ;
        RECT 75.000 17.100 75.400 17.200 ;
        RECT 74.200 16.800 75.400 17.100 ;
        RECT 72.300 16.200 72.600 16.800 ;
        RECT 75.000 16.400 75.400 16.800 ;
        RECT 75.800 16.200 76.100 17.500 ;
        RECT 71.500 15.900 72.000 16.200 ;
        RECT 72.300 15.900 73.000 16.200 ;
        RECT 67.800 14.800 68.200 15.600 ;
        RECT 68.600 14.200 68.900 15.900 ;
        RECT 71.700 14.200 72.000 15.900 ;
        RECT 72.600 15.800 73.000 15.900 ;
        RECT 75.800 15.800 76.200 16.200 ;
        RECT 76.600 16.100 77.000 16.200 ;
        RECT 77.400 16.100 77.800 19.900 ;
        RECT 79.500 19.200 79.900 19.900 ;
        RECT 79.500 18.800 80.200 19.200 ;
        RECT 79.500 16.300 79.900 18.800 ;
        RECT 76.600 15.800 77.800 16.100 ;
        RECT 79.000 15.900 79.900 16.300 ;
        RECT 80.600 16.200 81.000 19.900 ;
        RECT 81.300 16.200 81.700 16.300 ;
        RECT 80.600 15.900 81.700 16.200 ;
        RECT 82.800 16.200 83.600 19.900 ;
        RECT 84.600 16.200 85.000 16.300 ;
        RECT 85.400 16.200 85.800 19.900 ;
        RECT 86.600 16.800 87.000 17.200 ;
        RECT 86.600 16.200 86.900 16.800 ;
        RECT 87.300 16.200 87.700 19.900 ;
        RECT 82.800 15.900 83.800 16.200 ;
        RECT 84.600 15.900 85.800 16.200 ;
        RECT 86.200 15.900 86.900 16.200 ;
        RECT 87.200 15.900 87.700 16.200 ;
        RECT 72.600 14.800 73.000 15.200 ;
        RECT 74.200 14.800 75.400 15.200 ;
        RECT 72.600 14.200 72.900 14.800 ;
        RECT 75.800 14.200 76.100 15.800 ;
        RECT 68.600 13.800 69.000 14.200 ;
        RECT 70.200 14.100 70.600 14.200 ;
        RECT 69.400 13.800 71.000 14.100 ;
        RECT 71.700 13.800 73.000 14.200 ;
        RECT 75.300 14.100 76.100 14.200 ;
        RECT 75.200 13.900 76.100 14.100 ;
        RECT 68.600 12.200 68.900 13.800 ;
        RECT 69.400 13.200 69.700 13.800 ;
        RECT 70.600 13.600 71.000 13.800 ;
        RECT 69.400 12.400 69.800 13.200 ;
        RECT 70.300 13.100 72.100 13.300 ;
        RECT 72.600 13.100 72.900 13.800 ;
        RECT 70.200 13.000 72.200 13.100 ;
        RECT 68.600 11.100 69.000 12.200 ;
        RECT 70.200 11.100 70.600 13.000 ;
        RECT 71.800 11.100 72.200 13.000 ;
        RECT 72.600 11.100 73.000 13.100 ;
        RECT 75.200 11.100 75.600 13.900 ;
        RECT 76.600 12.400 77.000 13.200 ;
        RECT 77.400 11.100 77.800 15.800 ;
        RECT 79.100 14.200 79.400 15.900 ;
        RECT 81.400 15.600 81.700 15.900 ;
        RECT 81.400 15.300 83.100 15.600 ;
        RECT 82.700 15.200 83.100 15.300 ;
        RECT 83.500 15.200 83.800 15.900 ;
        RECT 86.200 15.800 86.600 15.900 ;
        RECT 83.500 15.100 84.200 15.200 ;
        RECT 86.200 15.100 86.600 15.200 ;
        RECT 81.600 14.900 82.000 15.000 ;
        RECT 83.500 14.900 86.600 15.100 ;
        RECT 81.600 14.600 82.900 14.900 ;
        RECT 82.600 14.300 82.900 14.600 ;
        RECT 83.300 14.800 86.600 14.900 ;
        RECT 83.300 14.600 83.800 14.800 ;
        RECT 79.000 13.800 79.400 14.200 ;
        RECT 80.600 14.100 81.400 14.200 ;
        RECT 80.600 13.800 82.300 14.100 ;
        RECT 82.600 13.900 83.000 14.300 ;
        RECT 79.100 12.100 79.400 13.800 ;
        RECT 82.000 13.600 82.300 13.800 ;
        RECT 81.300 13.400 81.700 13.500 ;
        RECT 79.000 11.100 79.400 12.100 ;
        RECT 80.600 13.100 81.700 13.400 ;
        RECT 82.000 13.300 83.000 13.600 ;
        RECT 82.200 13.200 83.000 13.300 ;
        RECT 80.600 11.100 81.000 13.100 ;
        RECT 83.300 12.900 83.600 14.600 ;
        RECT 87.200 14.200 87.500 15.900 ;
        RECT 87.800 14.400 88.200 15.200 ;
        RECT 84.000 13.800 84.400 14.200 ;
        RECT 85.000 13.800 85.800 14.200 ;
        RECT 86.200 13.800 87.500 14.200 ;
        RECT 88.600 14.100 89.000 14.200 ;
        RECT 88.200 13.800 89.000 14.100 ;
        RECT 84.000 13.600 84.300 13.800 ;
        RECT 83.900 13.200 84.300 13.600 ;
        RECT 84.600 13.400 85.000 13.500 ;
        RECT 84.600 13.100 85.800 13.400 ;
        RECT 86.300 13.100 86.600 13.800 ;
        RECT 88.200 13.600 88.600 13.800 ;
        RECT 89.400 13.400 89.800 14.200 ;
        RECT 87.100 13.100 88.900 13.300 ;
        RECT 82.800 11.100 83.600 12.900 ;
        RECT 85.400 11.100 85.800 13.100 ;
        RECT 86.200 11.100 86.600 13.100 ;
        RECT 87.000 13.000 89.000 13.100 ;
        RECT 87.000 11.100 87.400 13.000 ;
        RECT 88.600 11.100 89.000 13.000 ;
        RECT 90.200 11.100 90.600 19.900 ;
        RECT 91.000 16.200 91.400 19.900 ;
        RECT 92.600 16.200 93.000 19.900 ;
        RECT 91.000 15.900 93.000 16.200 ;
        RECT 93.400 15.900 93.800 19.900 ;
        RECT 94.600 16.800 95.000 17.200 ;
        RECT 94.600 16.200 94.900 16.800 ;
        RECT 95.300 16.200 95.700 19.900 ;
        RECT 94.200 15.900 94.900 16.200 ;
        RECT 95.200 15.900 95.700 16.200 ;
        RECT 97.400 15.900 97.800 19.900 ;
        RECT 99.000 17.900 99.400 19.900 ;
        RECT 91.400 15.200 91.800 15.400 ;
        RECT 93.400 15.200 93.700 15.900 ;
        RECT 94.200 15.800 94.600 15.900 ;
        RECT 91.000 14.900 91.800 15.200 ;
        RECT 92.600 14.900 93.800 15.200 ;
        RECT 91.000 14.800 91.400 14.900 ;
        RECT 91.000 14.200 91.300 14.800 ;
        RECT 91.000 13.800 91.400 14.200 ;
        RECT 91.800 13.800 92.200 14.600 ;
        RECT 92.600 13.100 92.900 14.900 ;
        RECT 93.400 14.800 93.800 14.900 ;
        RECT 95.200 14.200 95.500 15.900 ;
        RECT 97.400 15.200 97.700 15.900 ;
        RECT 99.000 15.800 99.300 17.900 ;
        RECT 103.500 16.300 103.900 19.900 ;
        RECT 105.900 17.200 106.300 19.900 ;
        RECT 105.400 16.800 106.300 17.200 ;
        RECT 106.600 16.800 107.400 17.200 ;
        RECT 103.000 15.900 103.900 16.300 ;
        RECT 105.900 16.200 106.300 16.800 ;
        RECT 106.700 16.200 107.000 16.800 ;
        RECT 109.100 16.200 109.500 19.900 ;
        RECT 109.800 16.800 110.200 17.200 ;
        RECT 109.900 16.200 110.200 16.800 ;
        RECT 105.900 15.900 106.400 16.200 ;
        RECT 106.700 15.900 107.400 16.200 ;
        RECT 109.100 15.900 109.600 16.200 ;
        RECT 109.900 15.900 110.600 16.200 ;
        RECT 112.300 15.900 113.300 19.900 ;
        RECT 115.300 17.200 115.700 19.900 ;
        RECT 115.300 16.800 116.200 17.200 ;
        RECT 115.300 16.300 115.700 16.800 ;
        RECT 115.300 15.900 116.200 16.300 ;
        RECT 117.400 15.900 117.800 19.900 ;
        RECT 119.000 17.900 119.400 19.900 ;
        RECT 98.100 15.500 99.300 15.800 ;
        RECT 95.800 14.400 96.200 15.200 ;
        RECT 97.400 15.100 97.800 15.200 ;
        RECT 96.600 14.800 97.800 15.100 ;
        RECT 94.200 13.800 95.500 14.200 ;
        RECT 96.600 14.200 96.900 14.800 ;
        RECT 96.600 14.100 97.000 14.200 ;
        RECT 96.200 13.800 97.000 14.100 ;
        RECT 93.400 13.100 93.800 13.200 ;
        RECT 94.300 13.100 94.600 13.800 ;
        RECT 96.200 13.600 96.600 13.800 ;
        RECT 95.100 13.100 96.900 13.300 ;
        RECT 97.400 13.100 97.700 14.800 ;
        RECT 98.100 13.800 98.400 15.500 ;
        RECT 99.000 14.800 99.400 15.200 ;
        RECT 101.400 15.100 101.800 15.200 ;
        RECT 103.100 15.100 103.400 15.900 ;
        RECT 101.400 14.800 103.400 15.100 ;
        RECT 103.800 15.100 104.200 15.600 ;
        RECT 104.600 15.100 105.000 15.200 ;
        RECT 103.800 14.800 105.000 15.100 ;
        RECT 99.000 14.400 99.300 14.800 ;
        RECT 98.800 14.100 99.300 14.400 ;
        RECT 98.800 14.000 99.200 14.100 ;
        RECT 99.800 13.800 100.200 14.600 ;
        RECT 103.100 14.200 103.400 14.800 ;
        RECT 105.400 14.400 105.800 15.200 ;
        RECT 106.100 14.200 106.400 15.900 ;
        RECT 107.000 15.800 107.400 15.900 ;
        RECT 107.000 15.100 107.400 15.200 ;
        RECT 108.600 15.100 109.000 15.200 ;
        RECT 107.000 14.800 109.000 15.100 ;
        RECT 108.600 14.400 109.000 14.800 ;
        RECT 109.300 14.200 109.600 15.900 ;
        RECT 110.200 15.800 110.600 15.900 ;
        RECT 110.200 15.200 110.500 15.800 ;
        RECT 110.200 14.800 110.600 15.200 ;
        RECT 103.000 13.800 103.400 14.200 ;
        RECT 104.600 14.100 105.000 14.200 ;
        RECT 104.600 13.800 105.400 14.100 ;
        RECT 106.100 13.800 107.400 14.200 ;
        RECT 107.800 14.100 108.200 14.200 ;
        RECT 107.800 13.800 108.600 14.100 ;
        RECT 109.300 13.800 110.600 14.200 ;
        RECT 111.000 13.800 111.400 14.600 ;
        RECT 111.800 14.400 112.200 15.200 ;
        RECT 112.700 14.200 113.000 15.900 ;
        RECT 113.400 14.400 113.800 15.200 ;
        RECT 115.000 14.800 115.400 15.600 ;
        RECT 115.800 14.200 116.100 15.900 ;
        RECT 117.400 15.200 117.700 15.900 ;
        RECT 119.000 15.800 119.300 17.900 ;
        RECT 119.800 17.100 120.200 17.200 ;
        RECT 120.900 17.100 121.300 19.900 ;
        RECT 119.800 16.800 121.300 17.100 ;
        RECT 120.900 16.300 121.300 16.800 ;
        RECT 120.900 15.900 121.800 16.300 ;
        RECT 118.100 15.500 119.300 15.800 ;
        RECT 117.400 14.800 117.800 15.200 ;
        RECT 112.600 14.100 113.000 14.200 ;
        RECT 114.200 14.100 114.600 14.200 ;
        RECT 111.800 13.800 113.000 14.100 ;
        RECT 113.800 13.800 114.600 14.100 ;
        RECT 115.800 13.800 116.200 14.200 ;
        RECT 98.000 13.700 98.400 13.800 ;
        RECT 98.000 13.500 99.500 13.700 ;
        RECT 98.000 13.400 100.100 13.500 ;
        RECT 99.200 13.200 100.100 13.400 ;
        RECT 99.800 13.100 100.100 13.200 ;
        RECT 92.600 11.100 93.000 13.100 ;
        RECT 93.400 12.800 94.600 13.100 ;
        RECT 93.300 12.400 93.700 12.800 ;
        RECT 94.200 11.100 94.600 12.800 ;
        RECT 95.000 13.000 97.000 13.100 ;
        RECT 95.000 11.100 95.400 13.000 ;
        RECT 96.600 11.100 97.000 13.000 ;
        RECT 97.400 12.600 98.100 13.100 ;
        RECT 97.700 11.100 98.100 12.600 ;
        RECT 99.800 11.100 100.200 13.100 ;
        RECT 102.200 12.400 102.600 13.200 ;
        RECT 103.100 12.100 103.400 13.800 ;
        RECT 105.000 13.600 105.400 13.800 ;
        RECT 104.700 13.100 106.500 13.300 ;
        RECT 107.000 13.100 107.300 13.800 ;
        RECT 108.200 13.600 108.600 13.800 ;
        RECT 107.900 13.100 109.700 13.300 ;
        RECT 110.200 13.100 110.500 13.800 ;
        RECT 111.800 13.100 112.100 13.800 ;
        RECT 113.800 13.600 114.200 13.800 ;
        RECT 112.700 13.100 114.500 13.300 ;
        RECT 103.000 11.100 103.400 12.100 ;
        RECT 104.600 13.000 106.600 13.100 ;
        RECT 104.600 11.100 105.000 13.000 ;
        RECT 106.200 11.100 106.600 13.000 ;
        RECT 107.000 11.100 107.400 13.100 ;
        RECT 107.800 13.000 109.800 13.100 ;
        RECT 107.800 11.100 108.200 13.000 ;
        RECT 109.400 11.100 109.800 13.000 ;
        RECT 110.200 11.100 110.600 13.100 ;
        RECT 111.000 11.400 111.400 13.100 ;
        RECT 111.800 11.700 112.200 13.100 ;
        RECT 112.600 13.000 114.600 13.100 ;
        RECT 112.600 11.400 113.000 13.000 ;
        RECT 111.000 11.100 113.000 11.400 ;
        RECT 114.200 11.100 114.600 13.000 ;
        RECT 115.800 12.100 116.100 13.800 ;
        RECT 116.600 12.400 117.000 13.200 ;
        RECT 117.400 13.100 117.700 14.800 ;
        RECT 118.100 13.800 118.400 15.500 ;
        RECT 119.000 14.800 119.400 15.200 ;
        RECT 120.600 14.800 121.000 15.600 ;
        RECT 119.000 14.400 119.300 14.800 ;
        RECT 118.800 14.100 119.300 14.400 ;
        RECT 119.800 14.100 120.200 14.600 ;
        RECT 121.400 14.200 121.700 15.900 ;
        RECT 120.600 14.100 121.000 14.200 ;
        RECT 118.800 14.000 119.200 14.100 ;
        RECT 119.800 13.800 121.000 14.100 ;
        RECT 121.400 13.800 121.800 14.200 ;
        RECT 118.000 13.700 118.400 13.800 ;
        RECT 118.000 13.500 119.500 13.700 ;
        RECT 118.000 13.400 120.100 13.500 ;
        RECT 119.200 13.200 120.100 13.400 ;
        RECT 119.800 13.100 120.100 13.200 ;
        RECT 117.400 12.600 118.100 13.100 ;
        RECT 117.700 12.200 118.100 12.600 ;
        RECT 115.800 11.100 116.200 12.100 ;
        RECT 117.400 11.800 118.100 12.200 ;
        RECT 117.700 11.100 118.100 11.800 ;
        RECT 119.800 11.100 120.200 13.100 ;
        RECT 121.400 12.100 121.700 13.800 ;
        RECT 122.200 13.100 122.600 13.200 ;
        RECT 123.000 13.100 123.400 19.900 ;
        RECT 125.900 19.200 126.300 19.900 ;
        RECT 125.900 18.800 126.600 19.200 ;
        RECT 125.900 16.300 126.300 18.800 ;
        RECT 125.400 15.900 126.300 16.300 ;
        RECT 125.500 14.200 125.800 15.900 ;
        RECT 126.200 15.100 126.600 15.600 ;
        RECT 127.000 15.100 127.400 15.200 ;
        RECT 126.200 14.800 127.400 15.100 ;
        RECT 123.800 14.100 124.200 14.200 ;
        RECT 125.400 14.100 125.800 14.200 ;
        RECT 123.800 13.800 125.800 14.100 ;
        RECT 126.200 14.100 126.600 14.200 ;
        RECT 127.000 14.100 127.400 14.200 ;
        RECT 126.200 13.800 127.400 14.100 ;
        RECT 123.800 13.400 124.200 13.800 ;
        RECT 122.200 12.800 123.400 13.100 ;
        RECT 122.200 12.400 122.600 12.800 ;
        RECT 121.400 11.100 121.800 12.100 ;
        RECT 123.000 11.100 123.400 12.800 ;
        RECT 124.600 12.400 125.000 13.200 ;
        RECT 125.500 12.100 125.800 13.800 ;
        RECT 127.000 13.400 127.400 13.800 ;
        RECT 125.400 11.100 125.800 12.100 ;
        RECT 127.800 11.100 128.200 19.900 ;
        RECT 129.900 16.200 130.300 19.900 ;
        RECT 132.600 17.900 133.000 19.900 ;
        RECT 132.700 17.800 133.000 17.900 ;
        RECT 134.200 17.900 134.600 19.900 ;
        RECT 134.200 17.800 134.500 17.900 ;
        RECT 132.700 17.500 134.500 17.800 ;
        RECT 133.400 16.400 133.800 17.200 ;
        RECT 134.200 16.200 134.500 17.500 ;
        RECT 136.300 16.300 136.700 19.900 ;
        RECT 129.900 15.900 130.400 16.200 ;
        RECT 128.600 15.100 129.000 15.200 ;
        RECT 129.400 15.100 129.800 15.200 ;
        RECT 128.600 14.800 129.800 15.100 ;
        RECT 129.400 14.400 129.800 14.800 ;
        RECT 130.100 14.200 130.400 15.900 ;
        RECT 131.800 15.400 132.200 16.200 ;
        RECT 134.200 15.800 134.600 16.200 ;
        RECT 135.800 15.900 136.700 16.300 ;
        RECT 138.700 16.200 139.700 19.900 ;
        RECT 141.400 16.900 141.800 19.900 ;
        RECT 141.500 16.600 141.800 16.900 ;
        RECT 143.000 19.600 145.000 19.900 ;
        RECT 143.000 16.900 143.400 19.600 ;
        RECT 143.800 16.900 144.200 19.300 ;
        RECT 144.600 17.000 145.000 19.600 ;
        RECT 145.500 19.600 147.300 19.900 ;
        RECT 145.500 19.500 145.800 19.600 ;
        RECT 143.000 16.600 143.300 16.900 ;
        RECT 141.500 16.300 143.300 16.600 ;
        RECT 143.900 16.700 144.200 16.900 ;
        RECT 145.400 16.700 145.800 19.500 ;
        RECT 147.000 19.500 147.300 19.600 ;
        RECT 143.900 16.500 145.800 16.700 ;
        RECT 146.200 16.500 146.600 19.300 ;
        RECT 147.000 16.500 147.400 19.500 ;
        RECT 143.900 16.400 145.700 16.500 ;
        RECT 138.200 15.900 139.700 16.200 ;
        RECT 146.200 16.200 146.500 16.500 ;
        RECT 148.100 16.300 148.500 19.900 ;
        RECT 146.200 16.100 146.600 16.200 ;
        RECT 132.600 14.800 133.800 15.200 ;
        RECT 134.200 14.200 134.500 15.800 ;
        RECT 135.000 15.100 135.400 15.200 ;
        RECT 135.900 15.100 136.200 15.900 ;
        RECT 138.200 15.800 139.400 15.900 ;
        RECT 135.000 14.800 136.200 15.100 ;
        RECT 136.600 14.800 137.000 15.600 ;
        RECT 135.900 14.200 136.200 14.800 ;
        RECT 128.600 14.100 129.000 14.200 ;
        RECT 128.600 13.800 129.400 14.100 ;
        RECT 130.100 13.800 131.400 14.200 ;
        RECT 133.700 14.100 134.500 14.200 ;
        RECT 135.000 14.100 135.400 14.200 ;
        RECT 133.600 13.800 135.400 14.100 ;
        RECT 135.800 13.800 136.200 14.200 ;
        RECT 137.400 13.800 137.800 14.600 ;
        RECT 138.200 14.400 138.600 15.200 ;
        RECT 139.100 14.200 139.400 15.800 ;
        RECT 144.900 15.800 146.600 16.100 ;
        RECT 148.100 15.900 149.000 16.300 ;
        RECT 139.800 14.400 140.200 15.200 ;
        RECT 143.800 14.800 144.600 15.200 ;
        RECT 139.000 14.100 139.400 14.200 ;
        RECT 140.600 14.100 141.000 14.200 ;
        RECT 138.200 13.800 139.400 14.100 ;
        RECT 140.200 13.800 141.000 14.100 ;
        RECT 142.200 14.100 142.600 14.200 ;
        RECT 143.000 14.100 143.800 14.200 ;
        RECT 142.200 13.800 143.800 14.100 ;
        RECT 129.000 13.600 129.400 13.800 ;
        RECT 128.700 13.100 130.500 13.300 ;
        RECT 131.000 13.200 131.300 13.800 ;
        RECT 128.600 13.000 130.600 13.100 ;
        RECT 128.600 11.100 129.000 13.000 ;
        RECT 130.200 11.100 130.600 13.000 ;
        RECT 131.000 11.100 131.400 13.200 ;
        RECT 133.600 11.100 134.000 13.800 ;
        RECT 135.000 12.400 135.400 13.200 ;
        RECT 135.900 12.100 136.200 13.800 ;
        RECT 138.200 13.100 138.500 13.800 ;
        RECT 140.200 13.600 140.600 13.800 ;
        RECT 139.100 13.100 140.900 13.300 ;
        RECT 135.800 11.100 136.200 12.100 ;
        RECT 137.400 11.400 137.800 13.100 ;
        RECT 138.200 11.700 138.600 13.100 ;
        RECT 139.000 13.000 141.000 13.100 ;
        RECT 139.000 11.400 139.400 13.000 ;
        RECT 137.400 11.100 139.400 11.400 ;
        RECT 140.600 11.100 141.000 13.000 ;
        RECT 142.200 12.800 143.400 13.200 ;
        RECT 144.900 12.500 145.200 15.800 ;
        RECT 147.800 14.800 148.200 15.600 ;
        RECT 148.600 15.200 148.900 15.900 ;
        RECT 148.600 14.800 149.000 15.200 ;
        RECT 143.200 12.200 145.200 12.500 ;
        RECT 143.200 12.100 143.500 12.200 ;
        RECT 143.000 11.800 143.500 12.100 ;
        RECT 144.600 12.100 145.200 12.200 ;
        RECT 148.600 14.200 148.900 14.800 ;
        RECT 148.600 13.800 149.000 14.200 ;
        RECT 148.600 12.100 148.900 13.800 ;
        RECT 143.000 11.100 143.400 11.800 ;
        RECT 144.600 11.100 145.000 12.100 ;
        RECT 148.600 11.100 149.000 12.100 ;
        RECT 0.600 7.900 1.000 9.900 ;
        RECT 2.800 8.100 3.600 9.900 ;
        RECT 0.600 7.600 1.700 7.900 ;
        RECT 2.200 7.700 3.000 7.800 ;
        RECT 1.300 7.500 1.700 7.600 ;
        RECT 2.000 7.400 3.000 7.700 ;
        RECT 2.000 7.200 2.300 7.400 ;
        RECT 0.600 6.900 2.300 7.200 ;
        RECT 0.600 6.800 1.400 6.900 ;
        RECT 2.600 6.700 3.000 7.100 ;
        RECT 2.600 6.400 2.900 6.700 ;
        RECT 1.600 6.100 2.900 6.400 ;
        RECT 3.300 6.400 3.600 8.100 ;
        RECT 5.400 7.900 5.800 9.900 ;
        RECT 3.900 7.400 4.300 7.800 ;
        RECT 4.600 7.600 5.800 7.900 ;
        RECT 6.200 7.900 6.600 9.900 ;
        RECT 8.400 9.200 9.200 9.900 ;
        RECT 7.800 8.800 9.200 9.200 ;
        RECT 8.400 8.100 9.200 8.800 ;
        RECT 6.200 7.600 7.500 7.900 ;
        RECT 4.600 7.500 5.000 7.600 ;
        RECT 7.100 7.500 7.500 7.600 ;
        RECT 7.800 7.400 8.600 7.800 ;
        RECT 4.000 7.200 4.300 7.400 ;
        RECT 4.000 6.800 4.400 7.200 ;
        RECT 5.000 6.800 5.800 7.200 ;
        RECT 6.200 7.100 7.000 7.200 ;
        RECT 8.900 7.100 9.200 8.100 ;
        RECT 11.000 7.900 11.400 9.900 ;
        RECT 12.600 9.100 13.000 9.200 ;
        RECT 14.200 9.100 14.600 9.900 ;
        RECT 15.800 9.200 16.200 9.900 ;
        RECT 12.600 8.800 14.600 9.100 ;
        RECT 15.700 8.900 16.200 9.200 ;
        RECT 15.700 8.800 16.000 8.900 ;
        RECT 9.500 7.400 9.900 7.800 ;
        RECT 10.200 7.600 11.400 7.900 ;
        RECT 14.000 8.500 16.000 8.800 ;
        RECT 10.200 7.500 10.600 7.600 ;
        RECT 6.200 7.000 7.300 7.100 ;
        RECT 6.200 6.800 8.400 7.000 ;
        RECT 7.000 6.700 8.400 6.800 ;
        RECT 8.000 6.600 8.400 6.700 ;
        RECT 8.700 6.800 9.200 7.100 ;
        RECT 9.600 7.200 9.900 7.400 ;
        RECT 9.600 6.800 10.000 7.200 ;
        RECT 10.600 7.100 11.400 7.200 ;
        RECT 11.800 7.100 12.200 7.200 ;
        RECT 10.600 6.800 12.200 7.100 ;
        RECT 3.300 6.200 3.800 6.400 ;
        RECT 8.700 6.200 9.000 6.800 ;
        RECT 3.300 6.100 4.200 6.200 ;
        RECT 1.600 6.000 2.000 6.100 ;
        RECT 3.500 5.800 4.200 6.100 ;
        RECT 7.300 6.100 7.700 6.200 ;
        RECT 7.300 5.800 8.100 6.100 ;
        RECT 8.600 5.800 9.000 6.200 ;
        RECT 2.700 5.700 3.100 5.800 ;
        RECT 1.400 5.400 3.100 5.700 ;
        RECT 1.400 5.100 1.700 5.400 ;
        RECT 3.500 5.100 3.800 5.800 ;
        RECT 7.700 5.700 8.100 5.800 ;
        RECT 8.700 5.100 9.000 5.800 ;
        RECT 14.000 5.200 14.300 8.500 ;
        RECT 16.100 7.800 17.000 8.200 ;
        RECT 18.200 7.900 18.600 9.900 ;
        RECT 20.400 8.100 21.200 9.900 ;
        RECT 18.200 7.600 19.400 7.900 ;
        RECT 19.000 7.500 19.400 7.600 ;
        RECT 19.700 7.400 20.100 7.800 ;
        RECT 19.700 7.200 20.000 7.400 ;
        RECT 15.400 7.100 16.200 7.200 ;
        RECT 17.400 7.100 17.800 7.200 ;
        RECT 15.400 6.800 17.800 7.100 ;
        RECT 18.200 6.800 19.000 7.200 ;
        RECT 19.600 6.800 20.000 7.200 ;
        RECT 20.400 6.400 20.700 8.100 ;
        RECT 23.000 7.900 23.400 9.900 ;
        RECT 21.000 7.700 21.800 7.800 ;
        RECT 21.000 7.400 22.000 7.700 ;
        RECT 22.300 7.600 23.400 7.900 ;
        RECT 23.800 7.800 24.200 8.600 ;
        RECT 22.300 7.500 22.700 7.600 ;
        RECT 21.700 7.200 22.000 7.400 ;
        RECT 21.000 6.700 21.400 7.100 ;
        RECT 21.700 6.900 23.400 7.200 ;
        RECT 22.600 6.800 23.400 6.900 ;
        RECT 20.200 6.200 20.700 6.400 ;
        RECT 14.600 5.800 15.400 6.200 ;
        RECT 19.800 6.100 20.700 6.200 ;
        RECT 21.100 6.400 21.400 6.700 ;
        RECT 21.100 6.100 22.400 6.400 ;
        RECT 19.800 5.800 20.500 6.100 ;
        RECT 22.000 6.000 22.400 6.100 ;
        RECT 0.600 4.800 1.700 5.100 ;
        RECT 0.600 1.100 1.000 4.800 ;
        RECT 1.300 4.700 1.700 4.800 ;
        RECT 2.800 4.800 3.800 5.100 ;
        RECT 4.600 4.800 5.800 5.100 ;
        RECT 2.800 1.100 3.600 4.800 ;
        RECT 4.600 4.700 5.000 4.800 ;
        RECT 5.400 1.100 5.800 4.800 ;
        RECT 6.200 4.800 7.500 5.100 ;
        RECT 6.200 1.100 6.600 4.800 ;
        RECT 7.100 4.700 7.500 4.800 ;
        RECT 8.400 1.100 9.200 5.100 ;
        RECT 10.200 4.800 11.400 5.100 ;
        RECT 12.600 4.900 14.300 5.200 ;
        RECT 20.200 5.100 20.500 5.800 ;
        RECT 20.900 5.700 21.300 5.800 ;
        RECT 20.900 5.400 22.600 5.700 ;
        RECT 22.300 5.100 22.600 5.400 ;
        RECT 12.600 4.800 13.000 4.900 ;
        RECT 10.200 4.700 10.600 4.800 ;
        RECT 11.000 1.100 11.400 4.800 ;
        RECT 12.700 4.500 13.000 4.800 ;
        RECT 18.200 4.800 19.400 5.100 ;
        RECT 20.200 4.800 21.200 5.100 ;
        RECT 13.500 4.500 15.300 4.600 ;
        RECT 11.800 1.500 12.200 4.500 ;
        RECT 12.600 1.700 13.000 4.500 ;
        RECT 13.400 4.300 15.300 4.500 ;
        RECT 11.900 1.400 12.200 1.500 ;
        RECT 13.400 1.500 13.800 4.300 ;
        RECT 15.000 4.100 15.300 4.300 ;
        RECT 15.900 4.400 17.700 4.700 ;
        RECT 15.900 4.100 16.200 4.400 ;
        RECT 13.400 1.400 13.700 1.500 ;
        RECT 11.900 1.100 13.700 1.400 ;
        RECT 14.200 1.400 14.600 4.000 ;
        RECT 15.000 1.700 15.400 4.100 ;
        RECT 15.800 1.400 16.200 4.100 ;
        RECT 14.200 1.100 16.200 1.400 ;
        RECT 17.400 4.100 17.700 4.400 ;
        RECT 17.400 1.100 17.800 4.100 ;
        RECT 18.200 1.100 18.600 4.800 ;
        RECT 19.000 4.700 19.400 4.800 ;
        RECT 20.400 1.100 21.200 4.800 ;
        RECT 22.300 4.800 23.400 5.100 ;
        RECT 22.300 4.700 22.700 4.800 ;
        RECT 23.000 1.100 23.400 4.800 ;
        RECT 24.600 1.100 25.000 9.900 ;
        RECT 25.400 7.900 25.800 9.900 ;
        RECT 26.200 8.000 26.600 9.900 ;
        RECT 27.800 8.000 28.200 9.900 ;
        RECT 26.200 7.900 28.200 8.000 ;
        RECT 28.600 7.900 29.000 9.900 ;
        RECT 30.800 8.100 31.600 9.900 ;
        RECT 25.500 7.200 25.800 7.900 ;
        RECT 26.300 7.700 28.100 7.900 ;
        RECT 28.600 7.600 29.900 7.900 ;
        RECT 29.500 7.500 29.900 7.600 ;
        RECT 30.200 7.400 31.000 7.800 ;
        RECT 27.400 7.200 27.800 7.400 ;
        RECT 25.400 6.800 26.700 7.200 ;
        RECT 27.400 6.900 28.200 7.200 ;
        RECT 27.800 6.800 28.200 6.900 ;
        RECT 28.600 7.100 29.400 7.200 ;
        RECT 31.300 7.100 31.600 8.100 ;
        RECT 33.400 7.900 33.800 9.900 ;
        RECT 35.800 9.200 36.200 9.900 ;
        RECT 35.800 8.900 36.300 9.200 ;
        RECT 36.000 8.800 36.300 8.900 ;
        RECT 37.400 8.900 37.800 9.900 ;
        RECT 43.000 8.900 43.400 9.900 ;
        RECT 44.600 9.200 45.000 9.900 ;
        RECT 37.400 8.800 38.000 8.900 ;
        RECT 36.000 8.500 38.000 8.800 ;
        RECT 31.900 7.400 32.300 7.800 ;
        RECT 32.600 7.600 33.800 7.900 ;
        RECT 35.000 7.800 35.900 8.200 ;
        RECT 32.600 7.500 33.000 7.600 ;
        RECT 28.600 7.000 29.700 7.100 ;
        RECT 28.600 6.800 30.800 7.000 ;
        RECT 25.400 5.100 25.800 5.200 ;
        RECT 26.400 5.100 26.700 6.800 ;
        RECT 29.400 6.700 30.800 6.800 ;
        RECT 30.400 6.600 30.800 6.700 ;
        RECT 31.100 6.800 31.600 7.100 ;
        RECT 32.000 7.200 32.300 7.400 ;
        RECT 37.700 7.200 38.000 8.500 ;
        RECT 32.000 6.800 32.400 7.200 ;
        RECT 33.000 6.800 33.800 7.200 ;
        RECT 35.800 6.800 36.600 7.200 ;
        RECT 37.400 6.800 38.000 7.200 ;
        RECT 27.000 5.800 27.400 6.600 ;
        RECT 31.100 6.200 31.400 6.800 ;
        RECT 29.700 6.100 30.100 6.200 ;
        RECT 29.700 5.800 30.500 6.100 ;
        RECT 31.000 5.800 31.400 6.200 ;
        RECT 36.600 5.800 37.400 6.200 ;
        RECT 30.100 5.700 30.500 5.800 ;
        RECT 31.100 5.200 31.400 5.800 ;
        RECT 30.200 5.100 31.400 5.200 ;
        RECT 37.700 5.200 38.000 6.800 ;
        RECT 42.800 8.800 43.400 8.900 ;
        RECT 44.500 8.900 45.000 9.200 ;
        RECT 44.500 8.800 44.800 8.900 ;
        RECT 42.800 8.500 44.800 8.800 ;
        RECT 42.800 5.200 43.100 8.500 ;
        RECT 44.900 7.800 45.800 8.200 ;
        RECT 47.000 8.000 47.400 9.900 ;
        RECT 48.600 8.000 49.000 9.900 ;
        RECT 47.000 7.900 49.000 8.000 ;
        RECT 49.400 7.900 49.800 9.900 ;
        RECT 52.100 8.200 52.500 9.900 ;
        RECT 52.100 7.900 53.000 8.200 ;
        RECT 44.200 6.800 45.000 7.200 ;
        RECT 45.400 7.100 45.700 7.800 ;
        RECT 47.100 7.700 48.900 7.900 ;
        RECT 47.400 7.200 47.800 7.400 ;
        RECT 49.400 7.200 49.700 7.900 ;
        RECT 47.000 7.100 47.800 7.200 ;
        RECT 45.400 6.900 47.800 7.100 ;
        RECT 45.400 6.800 47.400 6.900 ;
        RECT 48.500 6.800 49.800 7.200 ;
        RECT 43.400 6.100 44.200 6.200 ;
        RECT 47.800 6.100 48.200 6.600 ;
        RECT 43.400 5.800 48.200 6.100 ;
        RECT 25.400 4.800 26.100 5.100 ;
        RECT 26.400 4.800 26.900 5.100 ;
        RECT 25.800 4.200 26.100 4.800 ;
        RECT 25.800 3.800 26.200 4.200 ;
        RECT 26.500 1.100 26.900 4.800 ;
        RECT 28.600 4.800 29.900 5.100 ;
        RECT 30.200 4.800 31.600 5.100 ;
        RECT 28.600 1.100 29.000 4.800 ;
        RECT 29.500 4.700 29.900 4.800 ;
        RECT 30.800 1.100 31.600 4.800 ;
        RECT 32.600 4.800 33.800 5.100 ;
        RECT 37.700 4.900 39.400 5.200 ;
        RECT 32.600 4.700 33.000 4.800 ;
        RECT 33.400 1.100 33.800 4.800 ;
        RECT 39.000 4.800 39.400 4.900 ;
        RECT 39.800 5.100 40.200 5.200 ;
        RECT 41.400 5.100 43.100 5.200 ;
        RECT 48.500 5.100 48.800 6.800 ;
        RECT 49.400 6.100 49.800 6.200 ;
        RECT 52.600 6.100 53.000 7.900 ;
        RECT 54.200 7.600 54.600 9.900 ;
        RECT 55.800 8.200 56.200 9.900 ;
        RECT 58.700 9.200 59.100 9.900 ;
        RECT 58.200 8.800 59.100 9.200 ;
        RECT 58.700 8.200 59.100 8.800 ;
        RECT 55.800 7.900 56.300 8.200 ;
        RECT 53.400 6.800 53.800 7.600 ;
        RECT 54.200 7.300 55.500 7.600 ;
        RECT 49.400 5.800 53.000 6.100 ;
        RECT 49.400 5.200 49.700 5.800 ;
        RECT 49.400 5.100 49.800 5.200 ;
        RECT 39.800 4.900 43.100 5.100 ;
        RECT 39.800 4.800 41.800 4.900 ;
        RECT 34.300 4.400 36.100 4.700 ;
        RECT 34.300 4.100 34.600 4.400 ;
        RECT 34.200 1.100 34.600 4.100 ;
        RECT 35.800 4.100 36.100 4.400 ;
        RECT 36.700 4.500 38.500 4.600 ;
        RECT 39.000 4.500 39.300 4.800 ;
        RECT 41.500 4.500 41.800 4.800 ;
        RECT 48.300 4.800 48.800 5.100 ;
        RECT 49.100 4.800 49.800 5.100 ;
        RECT 42.300 4.500 44.100 4.600 ;
        RECT 36.700 4.300 38.600 4.500 ;
        RECT 36.700 4.100 37.000 4.300 ;
        RECT 35.800 1.400 36.200 4.100 ;
        RECT 36.600 1.700 37.000 4.100 ;
        RECT 37.400 1.400 37.800 4.000 ;
        RECT 38.200 1.500 38.600 4.300 ;
        RECT 39.000 1.700 39.400 4.500 ;
        RECT 35.800 1.100 37.800 1.400 ;
        RECT 38.300 1.400 38.600 1.500 ;
        RECT 39.800 1.500 40.200 4.500 ;
        RECT 40.600 1.500 41.000 4.500 ;
        RECT 41.400 1.700 41.800 4.500 ;
        RECT 42.200 4.300 44.100 4.500 ;
        RECT 39.800 1.400 40.100 1.500 ;
        RECT 38.300 1.100 40.100 1.400 ;
        RECT 40.700 1.400 41.000 1.500 ;
        RECT 42.200 1.500 42.600 4.300 ;
        RECT 43.800 4.100 44.100 4.300 ;
        RECT 44.700 4.400 46.500 4.700 ;
        RECT 44.700 4.100 45.000 4.400 ;
        RECT 42.200 1.400 42.500 1.500 ;
        RECT 40.700 1.100 42.500 1.400 ;
        RECT 43.000 1.400 43.400 4.000 ;
        RECT 43.800 1.700 44.200 4.100 ;
        RECT 44.600 1.400 45.000 4.100 ;
        RECT 43.000 1.100 45.000 1.400 ;
        RECT 46.200 4.100 46.500 4.400 ;
        RECT 46.200 1.100 46.600 4.100 ;
        RECT 48.300 1.100 48.700 4.800 ;
        RECT 49.100 4.200 49.400 4.800 ;
        RECT 49.000 3.800 49.400 4.200 ;
        RECT 52.600 1.100 53.000 5.800 ;
        RECT 55.200 6.500 55.500 7.300 ;
        RECT 56.000 7.200 56.300 7.900 ;
        RECT 58.200 7.900 59.100 8.200 ;
        RECT 55.800 7.100 56.300 7.200 ;
        RECT 56.600 7.100 57.000 7.200 ;
        RECT 55.800 6.800 57.000 7.100 ;
        RECT 55.200 6.100 55.700 6.500 ;
        RECT 55.200 5.100 55.500 6.100 ;
        RECT 56.000 5.100 56.300 6.800 ;
        RECT 54.200 4.800 55.500 5.100 ;
        RECT 54.200 1.100 54.600 4.800 ;
        RECT 55.800 4.600 56.300 5.100 ;
        RECT 55.800 1.100 56.200 4.600 ;
        RECT 58.200 1.100 58.600 7.900 ;
        RECT 59.800 7.600 60.200 9.900 ;
        RECT 61.400 8.200 61.800 9.900 ;
        RECT 64.300 9.200 64.700 9.900 ;
        RECT 64.300 8.800 65.000 9.200 ;
        RECT 66.200 8.800 66.600 9.900 ;
        RECT 64.300 8.200 64.700 8.800 ;
        RECT 61.400 7.900 61.900 8.200 ;
        RECT 59.800 7.300 61.100 7.600 ;
        RECT 60.800 6.500 61.100 7.300 ;
        RECT 61.600 7.200 61.900 7.900 ;
        RECT 63.800 7.900 64.700 8.200 ;
        RECT 61.400 7.100 61.900 7.200 ;
        RECT 63.000 7.100 63.400 7.600 ;
        RECT 61.400 6.800 63.400 7.100 ;
        RECT 60.800 6.100 61.300 6.500 ;
        RECT 60.800 5.100 61.100 6.100 ;
        RECT 61.600 5.100 61.900 6.800 ;
        RECT 59.800 4.800 61.100 5.100 ;
        RECT 59.800 1.100 60.200 4.800 ;
        RECT 61.400 4.600 61.900 5.100 ;
        RECT 61.400 1.100 61.800 4.600 ;
        RECT 63.800 1.100 64.200 7.900 ;
        RECT 66.300 7.200 66.600 8.800 ;
        RECT 66.200 6.800 66.600 7.200 ;
        RECT 66.300 5.100 66.600 6.800 ;
        RECT 68.600 8.100 69.000 9.900 ;
        RECT 70.200 8.900 70.600 9.900 ;
        RECT 69.400 8.100 69.800 8.600 ;
        RECT 68.600 7.800 69.800 8.100 ;
        RECT 66.200 4.700 67.100 5.100 ;
        RECT 66.700 1.100 67.100 4.700 ;
        RECT 68.600 1.100 69.000 7.800 ;
        RECT 70.300 7.200 70.600 8.900 ;
        RECT 70.200 6.800 70.600 7.200 ;
        RECT 70.300 6.200 70.600 6.800 ;
        RECT 70.200 5.800 70.600 6.200 ;
        RECT 70.300 5.100 70.600 5.800 ;
        RECT 71.000 6.100 71.400 6.200 ;
        RECT 71.800 6.100 72.200 9.900 ;
        RECT 74.200 8.900 74.600 9.900 ;
        RECT 74.300 7.200 74.600 8.900 ;
        RECT 75.800 8.000 76.200 9.900 ;
        RECT 77.400 8.000 77.800 9.900 ;
        RECT 75.800 7.900 77.800 8.000 ;
        RECT 75.900 7.700 77.700 7.900 ;
        RECT 78.200 7.800 78.600 9.900 ;
        RECT 79.000 8.000 79.400 9.900 ;
        RECT 80.600 8.000 81.000 9.900 ;
        RECT 79.000 7.900 81.000 8.000 ;
        RECT 81.400 7.900 81.800 9.900 ;
        RECT 83.000 8.800 83.400 9.900 ;
        RECT 76.200 7.200 76.600 7.400 ;
        RECT 78.200 7.200 78.500 7.800 ;
        RECT 79.100 7.700 80.900 7.900 ;
        RECT 79.400 7.200 79.800 7.400 ;
        RECT 81.400 7.200 81.700 7.900 ;
        RECT 82.200 7.800 82.600 8.600 ;
        RECT 83.100 7.200 83.400 8.800 ;
        RECT 84.600 7.800 85.000 8.600 ;
        RECT 74.200 6.800 74.600 7.200 ;
        RECT 75.800 6.900 76.600 7.200 ;
        RECT 75.800 6.800 76.200 6.900 ;
        RECT 77.300 6.800 78.600 7.200 ;
        RECT 79.000 6.900 79.800 7.200 ;
        RECT 79.000 6.800 79.400 6.900 ;
        RECT 80.500 6.800 81.800 7.200 ;
        RECT 83.000 6.800 83.400 7.200 ;
        RECT 71.000 5.800 72.200 6.100 ;
        RECT 73.400 6.100 73.800 6.200 ;
        RECT 74.300 6.100 74.600 6.800 ;
        RECT 73.400 5.800 74.600 6.100 ;
        RECT 71.000 5.400 71.400 5.800 ;
        RECT 70.200 4.700 71.100 5.100 ;
        RECT 70.700 1.100 71.100 4.700 ;
        RECT 71.800 1.100 72.200 5.800 ;
        RECT 74.300 5.100 74.600 5.800 ;
        RECT 77.300 5.100 77.600 6.800 ;
        RECT 79.800 5.800 80.200 6.600 ;
        RECT 80.500 5.200 80.800 6.800 ;
        RECT 78.200 5.100 78.600 5.200 ;
        RECT 74.200 4.700 75.100 5.100 ;
        RECT 74.700 1.100 75.100 4.700 ;
        RECT 77.100 4.800 77.600 5.100 ;
        RECT 77.900 4.800 78.600 5.100 ;
        RECT 79.800 4.800 80.800 5.200 ;
        RECT 81.400 5.100 81.800 5.200 ;
        RECT 83.100 5.100 83.400 6.800 ;
        RECT 85.400 7.100 85.800 9.900 ;
        RECT 87.000 8.800 87.400 9.900 ;
        RECT 86.200 7.800 86.600 8.200 ;
        RECT 86.200 7.100 86.500 7.800 ;
        RECT 85.400 6.800 86.500 7.100 ;
        RECT 87.000 7.200 87.300 8.800 ;
        RECT 87.800 8.100 88.200 8.600 ;
        RECT 88.600 8.100 89.000 9.900 ;
        RECT 87.800 7.800 89.000 8.100 ;
        RECT 89.400 8.000 89.800 9.900 ;
        RECT 91.000 8.000 91.400 9.900 ;
        RECT 89.400 7.900 91.400 8.000 ;
        RECT 91.800 7.900 92.200 9.900 ;
        RECT 92.600 8.000 93.000 9.900 ;
        RECT 94.200 8.000 94.600 9.900 ;
        RECT 92.600 7.900 94.600 8.000 ;
        RECT 95.000 9.600 97.000 9.900 ;
        RECT 95.000 7.900 95.400 9.600 ;
        RECT 95.800 7.900 96.200 9.300 ;
        RECT 96.600 8.000 97.000 9.600 ;
        RECT 98.200 8.000 98.600 9.900 ;
        RECT 96.600 7.900 98.600 8.000 ;
        RECT 100.600 8.000 101.000 9.900 ;
        RECT 102.200 8.000 102.600 9.900 ;
        RECT 100.600 7.900 102.600 8.000 ;
        RECT 103.000 7.900 103.400 9.900 ;
        RECT 88.700 7.200 89.000 7.800 ;
        RECT 89.500 7.700 91.300 7.900 ;
        RECT 90.600 7.200 91.000 7.400 ;
        RECT 91.900 7.200 92.200 7.900 ;
        RECT 92.700 7.700 94.500 7.900 ;
        RECT 93.800 7.200 94.200 7.400 ;
        RECT 95.800 7.200 96.100 7.900 ;
        RECT 96.700 7.700 98.500 7.900 ;
        RECT 100.700 7.700 102.500 7.900 ;
        RECT 97.800 7.200 98.200 7.400 ;
        RECT 101.000 7.200 101.400 7.400 ;
        RECT 103.000 7.200 103.300 7.900 ;
        RECT 87.000 6.800 87.400 7.200 ;
        RECT 88.600 6.800 89.900 7.200 ;
        RECT 90.600 6.900 91.400 7.200 ;
        RECT 91.000 6.800 91.400 6.900 ;
        RECT 91.800 6.800 93.100 7.200 ;
        RECT 93.800 6.900 94.600 7.200 ;
        RECT 94.200 6.800 94.600 6.900 ;
        RECT 83.800 6.100 84.200 6.200 ;
        RECT 84.600 6.100 85.000 6.200 ;
        RECT 83.800 5.800 85.000 6.100 ;
        RECT 83.800 5.400 84.200 5.800 ;
        RECT 81.100 4.800 81.800 5.100 ;
        RECT 77.100 1.100 77.500 4.800 ;
        RECT 77.900 4.200 78.200 4.800 ;
        RECT 77.800 3.800 78.200 4.200 ;
        RECT 80.300 1.100 80.700 4.800 ;
        RECT 81.100 4.200 81.400 4.800 ;
        RECT 83.000 4.700 83.900 5.100 ;
        RECT 81.000 3.800 81.400 4.200 ;
        RECT 83.500 1.100 83.900 4.700 ;
        RECT 85.400 1.100 85.800 6.800 ;
        RECT 86.200 5.400 86.600 6.200 ;
        RECT 87.000 5.100 87.300 6.800 ;
        RECT 89.600 5.100 89.900 6.800 ;
        RECT 90.200 6.100 90.600 6.600 ;
        RECT 90.200 5.800 92.100 6.100 ;
        RECT 91.800 5.200 92.100 5.800 ;
        RECT 91.800 5.100 92.200 5.200 ;
        RECT 92.800 5.100 93.100 6.800 ;
        RECT 93.400 5.800 93.800 6.600 ;
        RECT 95.000 6.400 95.400 7.200 ;
        RECT 95.800 6.900 97.000 7.200 ;
        RECT 97.800 6.900 98.600 7.200 ;
        RECT 96.600 6.800 97.000 6.900 ;
        RECT 98.200 6.800 98.600 6.900 ;
        RECT 100.600 6.900 101.400 7.200 ;
        RECT 100.600 6.800 101.000 6.900 ;
        RECT 102.100 6.800 103.400 7.200 ;
        RECT 103.800 7.100 104.200 9.900 ;
        RECT 104.600 7.800 105.000 8.600 ;
        RECT 105.400 8.000 105.800 9.900 ;
        RECT 107.000 8.000 107.400 9.900 ;
        RECT 105.400 7.900 107.400 8.000 ;
        RECT 107.800 8.100 108.200 9.900 ;
        RECT 109.400 8.800 109.800 9.900 ;
        RECT 108.600 8.100 109.000 8.600 ;
        RECT 105.500 7.700 107.300 7.900 ;
        RECT 107.800 7.800 109.000 8.100 ;
        RECT 105.800 7.200 106.200 7.400 ;
        RECT 107.800 7.200 108.100 7.800 ;
        RECT 109.500 7.200 109.800 8.800 ;
        RECT 111.000 7.800 111.400 8.600 ;
        RECT 105.400 7.100 106.200 7.200 ;
        RECT 103.800 6.900 106.200 7.100 ;
        RECT 103.800 6.800 105.800 6.900 ;
        RECT 106.900 6.800 108.200 7.200 ;
        RECT 109.400 6.800 109.800 7.200 ;
        RECT 95.800 5.800 96.200 6.600 ;
        RECT 96.700 5.100 97.000 6.800 ;
        RECT 97.400 6.100 97.800 6.600 ;
        RECT 99.000 6.100 99.400 6.200 ;
        RECT 97.400 5.800 99.400 6.100 ;
        RECT 101.400 5.800 101.800 6.600 ;
        RECT 102.100 5.100 102.400 6.800 ;
        RECT 103.000 6.100 103.400 6.200 ;
        RECT 103.800 6.100 104.200 6.800 ;
        RECT 103.000 5.800 104.200 6.100 ;
        RECT 106.200 5.800 106.600 6.600 ;
        RECT 86.500 4.700 87.400 5.100 ;
        RECT 89.600 4.800 90.100 5.100 ;
        RECT 91.800 4.800 92.500 5.100 ;
        RECT 92.800 4.800 93.300 5.100 ;
        RECT 86.500 1.100 86.900 4.700 ;
        RECT 89.700 1.100 90.100 4.800 ;
        RECT 92.200 4.200 92.500 4.800 ;
        RECT 92.200 3.800 92.600 4.200 ;
        RECT 92.900 1.100 93.300 4.800 ;
        RECT 96.300 1.100 97.300 5.100 ;
        RECT 101.900 4.800 102.400 5.100 ;
        RECT 101.900 1.100 102.300 4.800 ;
        RECT 103.800 1.100 104.200 5.800 ;
        RECT 106.900 5.100 107.200 6.800 ;
        RECT 107.800 5.100 108.200 5.200 ;
        RECT 109.500 5.100 109.800 6.800 ;
        RECT 110.200 5.400 110.600 6.200 ;
        RECT 111.800 6.100 112.200 9.900 ;
        RECT 112.600 8.000 113.000 9.900 ;
        RECT 114.200 9.600 116.200 9.900 ;
        RECT 114.200 8.000 114.600 9.600 ;
        RECT 112.600 7.900 114.600 8.000 ;
        RECT 112.700 7.700 114.500 7.900 ;
        RECT 115.000 7.800 115.400 9.300 ;
        RECT 115.800 7.900 116.200 9.600 ;
        RECT 117.400 8.900 117.800 9.900 ;
        RECT 116.600 7.800 117.000 8.600 ;
        RECT 117.500 7.800 117.800 8.900 ;
        RECT 119.000 7.900 119.400 9.900 ;
        RECT 119.800 7.900 120.200 9.900 ;
        RECT 120.600 8.000 121.000 9.900 ;
        RECT 122.200 8.000 122.600 9.900 ;
        RECT 123.800 8.900 124.200 9.900 ;
        RECT 120.600 7.900 122.600 8.000 ;
        RECT 113.000 7.200 113.400 7.400 ;
        RECT 115.100 7.200 115.400 7.800 ;
        RECT 117.500 7.500 118.700 7.800 ;
        RECT 112.600 6.900 113.400 7.200 ;
        RECT 114.200 6.900 115.400 7.200 ;
        RECT 112.600 6.800 113.000 6.900 ;
        RECT 114.200 6.800 114.600 6.900 ;
        RECT 113.400 6.100 113.800 6.600 ;
        RECT 111.800 5.800 113.800 6.100 ;
        RECT 106.700 4.800 107.200 5.100 ;
        RECT 107.500 4.800 108.200 5.100 ;
        RECT 106.700 1.100 107.100 4.800 ;
        RECT 107.500 4.200 107.800 4.800 ;
        RECT 109.400 4.700 110.300 5.100 ;
        RECT 107.400 3.800 107.800 4.200 ;
        RECT 109.900 1.100 110.300 4.700 ;
        RECT 111.800 1.100 112.200 5.800 ;
        RECT 114.200 5.100 114.500 6.800 ;
        RECT 115.000 5.800 115.400 6.600 ;
        RECT 115.800 6.400 116.200 7.200 ;
        RECT 117.400 6.800 117.900 7.200 ;
        RECT 117.600 6.400 118.000 6.800 ;
        RECT 118.400 6.000 118.700 7.500 ;
        RECT 119.100 6.200 119.400 7.900 ;
        RECT 119.900 7.200 120.200 7.900 ;
        RECT 120.700 7.700 122.500 7.900 ;
        RECT 121.800 7.200 122.200 7.400 ;
        RECT 123.900 7.200 124.200 8.900 ;
        RECT 126.700 8.200 127.100 9.900 ;
        RECT 118.300 5.700 118.700 6.000 ;
        RECT 119.000 5.800 119.400 6.200 ;
        RECT 119.800 6.800 121.100 7.200 ;
        RECT 121.800 6.900 122.600 7.200 ;
        RECT 122.200 6.800 122.600 6.900 ;
        RECT 123.000 7.100 123.400 7.200 ;
        RECT 123.800 7.100 124.200 7.200 ;
        RECT 123.000 6.800 124.200 7.100 ;
        RECT 119.800 6.200 120.100 6.800 ;
        RECT 119.800 5.800 120.200 6.200 ;
        RECT 116.600 5.600 118.700 5.700 ;
        RECT 116.600 5.400 118.600 5.600 ;
        RECT 113.900 1.100 114.900 5.100 ;
        RECT 116.600 1.100 117.000 5.400 ;
        RECT 119.100 5.100 119.400 5.800 ;
        RECT 118.700 4.800 119.400 5.100 ;
        RECT 120.800 5.100 121.100 6.800 ;
        RECT 121.400 5.800 121.800 6.600 ;
        RECT 123.900 5.100 124.200 6.800 ;
        RECT 126.200 8.100 127.100 8.200 ;
        RECT 127.800 8.100 128.200 8.600 ;
        RECT 126.200 7.800 128.200 8.100 ;
        RECT 120.800 4.800 121.300 5.100 ;
        RECT 118.700 1.100 119.100 4.800 ;
        RECT 120.900 1.100 121.300 4.800 ;
        RECT 123.800 4.700 124.700 5.100 ;
        RECT 124.300 1.100 124.700 4.700 ;
        RECT 126.200 1.100 126.600 7.800 ;
        RECT 128.600 6.100 129.000 9.900 ;
        RECT 129.400 8.000 129.800 9.900 ;
        RECT 131.000 8.000 131.400 9.900 ;
        RECT 129.400 7.900 131.400 8.000 ;
        RECT 131.800 7.900 132.200 9.900 ;
        RECT 133.400 8.900 133.800 9.900 ;
        RECT 129.500 7.700 131.300 7.900 ;
        RECT 129.800 7.200 130.200 7.400 ;
        RECT 131.800 7.200 132.100 7.900 ;
        RECT 133.400 7.200 133.700 8.900 ;
        RECT 134.200 7.800 134.600 8.600 ;
        RECT 129.400 6.900 130.200 7.200 ;
        RECT 130.900 7.100 132.200 7.200 ;
        RECT 132.600 7.100 133.000 7.200 ;
        RECT 129.400 6.800 129.800 6.900 ;
        RECT 130.900 6.800 133.000 7.100 ;
        RECT 133.400 7.100 133.800 7.200 ;
        RECT 135.000 7.100 135.400 7.600 ;
        RECT 133.400 6.800 135.400 7.100 ;
        RECT 135.800 7.100 136.200 9.900 ;
        RECT 137.400 8.900 137.800 9.900 ;
        RECT 136.600 7.800 137.000 8.600 ;
        RECT 137.500 7.800 137.800 8.900 ;
        RECT 139.000 7.900 139.400 9.900 ;
        RECT 137.500 7.500 138.700 7.800 ;
        RECT 137.400 7.100 137.900 7.200 ;
        RECT 135.800 6.800 137.900 7.100 ;
        RECT 130.200 6.100 130.600 6.600 ;
        RECT 128.600 5.800 130.600 6.100 ;
        RECT 128.600 1.100 129.000 5.800 ;
        RECT 130.900 5.100 131.200 6.800 ;
        RECT 132.600 5.400 133.000 6.200 ;
        RECT 131.800 5.100 132.200 5.200 ;
        RECT 133.400 5.100 133.700 6.800 ;
        RECT 130.700 4.800 131.200 5.100 ;
        RECT 131.500 4.800 132.200 5.100 ;
        RECT 130.700 1.100 131.100 4.800 ;
        RECT 131.500 4.200 131.800 4.800 ;
        RECT 131.400 3.800 131.800 4.200 ;
        RECT 132.900 4.700 133.800 5.100 ;
        RECT 132.900 1.100 133.300 4.700 ;
        RECT 135.800 1.100 136.200 6.800 ;
        RECT 137.600 6.400 138.000 6.800 ;
        RECT 138.400 6.000 138.700 7.500 ;
        RECT 139.100 7.100 139.400 7.900 ;
        RECT 141.400 7.900 141.800 9.900 ;
        RECT 142.100 8.200 142.500 8.600 ;
        RECT 140.600 7.100 141.000 7.200 ;
        RECT 139.000 6.800 141.000 7.100 ;
        RECT 139.100 6.200 139.400 6.800 ;
        RECT 140.600 6.400 141.000 6.800 ;
        RECT 138.300 5.700 138.700 6.000 ;
        RECT 139.000 5.800 139.400 6.200 ;
        RECT 139.800 6.100 140.200 6.200 ;
        RECT 141.400 6.100 141.700 7.900 ;
        RECT 142.200 7.800 142.600 8.200 ;
        RECT 144.600 7.900 145.000 9.900 ;
        RECT 145.300 8.200 145.700 8.600 ;
        RECT 143.800 6.400 144.200 7.200 ;
        RECT 142.200 6.100 142.600 6.200 ;
        RECT 139.800 5.800 140.600 6.100 ;
        RECT 141.400 5.800 142.600 6.100 ;
        RECT 143.000 6.100 143.400 6.200 ;
        RECT 144.600 6.100 144.900 7.900 ;
        RECT 145.400 7.800 145.800 8.200 ;
        RECT 146.200 8.000 146.600 9.900 ;
        RECT 147.800 8.000 148.200 9.900 ;
        RECT 146.200 7.900 148.200 8.000 ;
        RECT 148.600 7.900 149.000 9.900 ;
        RECT 146.300 7.700 148.100 7.900 ;
        RECT 146.600 7.200 147.000 7.400 ;
        RECT 148.600 7.200 148.900 7.900 ;
        RECT 146.200 6.900 147.000 7.200 ;
        RECT 146.200 6.800 146.600 6.900 ;
        RECT 147.700 6.800 149.000 7.200 ;
        RECT 145.400 6.100 145.800 6.200 ;
        RECT 143.000 5.800 143.800 6.100 ;
        RECT 144.600 5.800 145.800 6.100 ;
        RECT 147.000 5.800 147.400 6.600 ;
        RECT 136.600 5.600 138.700 5.700 ;
        RECT 136.600 5.400 138.600 5.600 ;
        RECT 136.600 1.100 137.000 5.400 ;
        RECT 139.100 5.100 139.400 5.800 ;
        RECT 140.200 5.600 140.600 5.800 ;
        RECT 142.200 5.100 142.500 5.800 ;
        RECT 143.400 5.600 143.800 5.800 ;
        RECT 145.400 5.100 145.700 5.800 ;
        RECT 147.700 5.100 148.000 6.800 ;
        RECT 148.600 5.100 149.000 5.200 ;
        RECT 149.400 5.100 149.800 5.200 ;
        RECT 138.700 4.800 139.400 5.100 ;
        RECT 139.800 4.800 141.800 5.100 ;
        RECT 138.700 1.100 139.100 4.800 ;
        RECT 139.800 1.100 140.200 4.800 ;
        RECT 141.400 1.100 141.800 4.800 ;
        RECT 142.200 1.100 142.600 5.100 ;
        RECT 143.000 4.800 145.000 5.100 ;
        RECT 143.000 1.100 143.400 4.800 ;
        RECT 144.600 1.100 145.000 4.800 ;
        RECT 145.400 1.100 145.800 5.100 ;
        RECT 147.500 4.800 148.000 5.100 ;
        RECT 148.300 4.800 149.800 5.100 ;
        RECT 147.500 1.100 147.900 4.800 ;
        RECT 148.300 4.200 148.600 4.800 ;
        RECT 148.200 3.800 148.600 4.200 ;
      LAYER via1 ;
        RECT 4.600 126.800 5.000 127.200 ;
        RECT 7.000 126.800 7.400 127.200 ;
        RECT 2.200 125.800 2.600 126.200 ;
        RECT 8.600 126.800 9.000 127.200 ;
        RECT 15.800 126.800 16.200 127.200 ;
        RECT 7.000 121.800 7.400 122.200 ;
        RECT 18.200 125.800 18.600 126.200 ;
        RECT 15.800 124.800 16.200 125.200 ;
        RECT 26.200 125.800 26.600 126.200 ;
        RECT 29.400 125.800 29.800 126.200 ;
        RECT 30.200 125.800 30.600 126.200 ;
        RECT 23.800 124.800 24.200 125.200 ;
        RECT 47.000 128.800 47.400 129.200 ;
        RECT 46.200 126.800 46.600 127.200 ;
        RECT 22.200 123.800 22.600 124.200 ;
        RECT 18.200 121.800 18.600 122.200 ;
        RECT 36.600 124.900 37.000 125.300 ;
        RECT 40.600 125.800 41.000 126.200 ;
        RECT 61.400 127.800 61.800 128.200 ;
        RECT 40.600 123.800 41.000 124.200 ;
        RECT 44.600 124.800 45.000 125.200 ;
        RECT 55.000 125.800 55.400 126.200 ;
        RECT 65.400 126.800 65.800 127.200 ;
        RECT 59.800 125.800 60.200 126.200 ;
        RECT 55.000 121.800 55.400 122.200 ;
        RECT 65.400 124.800 65.800 125.200 ;
        RECT 74.200 125.800 74.600 126.200 ;
        RECT 71.000 124.800 71.400 125.200 ;
        RECT 74.200 121.800 74.600 122.200 ;
        RECT 87.000 126.500 87.400 126.900 ;
        RECT 81.400 125.800 81.800 126.200 ;
        RECT 91.800 126.300 92.200 126.700 ;
        RECT 84.600 125.800 85.000 126.200 ;
        RECT 87.800 124.400 88.200 124.800 ;
        RECT 90.200 123.800 90.600 124.200 ;
        RECT 81.400 121.800 81.800 122.200 ;
        RECT 88.600 123.100 89.000 123.500 ;
        RECT 87.000 122.100 87.400 122.500 ;
        RECT 87.800 122.100 88.200 122.500 ;
        RECT 90.200 123.100 90.600 123.500 ;
        RECT 91.800 123.100 92.200 123.500 ;
        RECT 92.600 122.100 93.000 122.500 ;
        RECT 93.400 122.100 93.800 122.500 ;
        RECT 94.200 122.100 94.600 122.500 ;
        RECT 106.200 126.500 106.600 126.900 ;
        RECT 111.000 126.300 111.400 126.700 ;
        RECT 103.800 125.800 104.200 126.200 ;
        RECT 107.000 124.400 107.400 124.800 ;
        RECT 109.400 123.800 109.800 124.200 ;
        RECT 99.000 121.800 99.400 122.200 ;
        RECT 107.800 123.100 108.200 123.500 ;
        RECT 106.200 122.100 106.600 122.500 ;
        RECT 107.000 122.100 107.400 122.500 ;
        RECT 109.400 123.100 109.800 123.500 ;
        RECT 111.000 123.100 111.400 123.500 ;
        RECT 111.800 122.100 112.200 122.500 ;
        RECT 112.600 122.100 113.000 122.500 ;
        RECT 113.400 122.100 113.800 122.500 ;
        RECT 118.200 121.800 118.600 122.200 ;
        RECT 125.400 126.500 125.800 126.900 ;
        RECT 130.200 126.300 130.600 126.700 ;
        RECT 138.200 127.800 138.600 128.200 ;
        RECT 123.000 125.800 123.400 126.200 ;
        RECT 124.600 125.800 125.000 126.200 ;
        RECT 126.200 124.400 126.600 124.800 ;
        RECT 128.600 123.800 129.000 124.200 ;
        RECT 119.800 121.800 120.200 122.200 ;
        RECT 127.000 123.100 127.400 123.500 ;
        RECT 125.400 122.100 125.800 122.500 ;
        RECT 126.200 122.100 126.600 122.500 ;
        RECT 128.600 123.100 129.000 123.500 ;
        RECT 130.200 123.100 130.600 123.500 ;
        RECT 131.000 122.100 131.400 122.500 ;
        RECT 131.800 122.100 132.200 122.500 ;
        RECT 132.600 122.100 133.000 122.500 ;
        RECT 147.800 124.800 148.200 125.200 ;
        RECT 147.000 121.800 147.400 122.200 ;
        RECT 148.600 121.800 149.000 122.200 ;
        RECT 2.200 118.800 2.600 119.200 ;
        RECT 1.400 116.800 1.800 117.200 ;
        RECT 4.600 116.800 5.000 117.200 ;
        RECT 9.400 118.800 9.800 119.200 ;
        RECT 3.000 115.800 3.400 116.200 ;
        RECT 6.200 115.800 6.600 116.200 ;
        RECT 2.200 114.800 2.600 115.200 ;
        RECT 5.400 114.800 5.800 115.200 ;
        RECT 12.600 116.800 13.000 117.200 ;
        RECT 11.800 115.800 12.200 116.200 ;
        RECT 11.000 114.800 11.400 115.200 ;
        RECT 8.600 112.800 9.000 113.200 ;
        RECT 7.800 111.800 8.200 112.200 ;
        RECT 17.400 118.800 17.800 119.200 ;
        RECT 16.600 114.800 17.000 115.200 ;
        RECT 25.400 116.800 25.800 117.200 ;
        RECT 14.200 113.800 14.600 114.200 ;
        RECT 20.600 113.800 21.000 114.200 ;
        RECT 21.400 113.800 21.800 114.200 ;
        RECT 18.200 112.800 18.600 113.200 ;
        RECT 23.000 113.800 23.400 114.200 ;
        RECT 31.800 118.800 32.200 119.200 ;
        RECT 38.200 118.800 38.600 119.200 ;
        RECT 40.600 118.800 41.000 119.200 ;
        RECT 33.400 116.800 33.800 117.200 ;
        RECT 37.400 116.800 37.800 117.200 ;
        RECT 35.000 115.800 35.400 116.200 ;
        RECT 35.800 115.800 36.200 116.200 ;
        RECT 44.600 118.800 45.000 119.200 ;
        RECT 43.800 116.800 44.200 117.200 ;
        RECT 34.200 114.800 34.600 115.200 ;
        RECT 42.200 115.800 42.600 116.200 ;
        RECT 40.600 114.800 41.000 115.200 ;
        RECT 33.400 113.800 33.800 114.200 ;
        RECT 41.400 113.800 41.800 114.200 ;
        RECT 46.200 111.800 46.600 112.200 ;
        RECT 55.000 118.800 55.400 119.200 ;
        RECT 51.800 113.800 52.200 114.200 ;
        RECT 51.000 112.800 51.400 113.200 ;
        RECT 59.000 118.800 59.400 119.200 ;
        RECT 57.400 113.800 57.800 114.200 ;
        RECT 50.200 111.800 50.600 112.200 ;
        RECT 64.600 118.800 65.000 119.200 ;
        RECT 69.400 116.800 69.800 117.200 ;
        RECT 75.800 118.800 76.200 119.200 ;
        RECT 67.800 115.800 68.200 116.200 ;
        RECT 75.000 116.800 75.400 117.200 ;
        RECT 56.600 112.800 57.000 113.200 ;
        RECT 63.800 113.800 64.200 114.200 ;
        RECT 63.000 112.800 63.400 113.200 ;
        RECT 71.000 114.800 71.400 115.200 ;
        RECT 71.800 114.800 72.200 115.200 ;
        RECT 76.600 115.800 77.000 116.200 ;
        RECT 75.800 114.800 76.200 115.200 ;
        RECT 80.600 114.800 81.000 115.200 ;
        RECT 91.000 117.500 91.400 117.900 ;
        RECT 89.400 116.800 89.800 117.200 ;
        RECT 91.800 116.200 92.200 116.600 ;
        RECT 102.200 116.800 102.600 117.200 ;
        RECT 86.200 114.100 86.600 114.500 ;
        RECT 91.000 114.300 91.400 114.700 ;
        RECT 77.400 112.800 77.800 113.200 ;
        RECT 88.600 113.800 89.000 114.200 ;
        RECT 86.200 112.100 86.600 112.500 ;
        RECT 87.000 112.100 87.400 112.500 ;
        RECT 87.800 112.100 88.200 112.500 ;
        RECT 89.400 112.100 89.800 112.500 ;
        RECT 91.000 112.100 91.400 112.500 ;
        RECT 91.800 112.100 92.200 112.500 ;
        RECT 92.600 112.100 93.000 112.500 ;
        RECT 93.400 112.100 93.800 112.500 ;
        RECT 106.200 118.800 106.600 119.200 ;
        RECT 110.200 116.800 110.600 117.200 ;
        RECT 105.400 113.800 105.800 114.200 ;
        RECT 98.200 111.800 98.600 112.200 ;
        RECT 103.000 112.800 103.400 113.200 ;
        RECT 111.800 115.800 112.200 116.200 ;
        RECT 111.000 114.800 111.400 115.200 ;
        RECT 111.000 111.800 111.400 112.200 ;
        RECT 116.600 118.800 117.000 119.200 ;
        RECT 113.400 112.800 113.800 113.200 ;
        RECT 131.000 117.500 131.400 117.900 ;
        RECT 129.400 116.800 129.800 117.200 ;
        RECT 131.800 116.200 132.200 116.600 ;
        RECT 126.200 114.100 126.600 114.500 ;
        RECT 131.000 114.300 131.400 114.700 ;
        RECT 128.600 113.800 129.000 114.200 ;
        RECT 139.000 113.800 139.400 114.200 ;
        RECT 126.200 112.100 126.600 112.500 ;
        RECT 127.000 112.100 127.400 112.500 ;
        RECT 127.800 112.100 128.200 112.500 ;
        RECT 129.400 112.100 129.800 112.500 ;
        RECT 131.000 112.100 131.400 112.500 ;
        RECT 131.800 112.100 132.200 112.500 ;
        RECT 132.600 112.100 133.000 112.500 ;
        RECT 133.400 112.100 133.800 112.500 ;
        RECT 143.800 114.800 144.200 115.200 ;
        RECT 146.200 114.800 146.600 115.200 ;
        RECT 140.600 112.800 141.000 113.200 ;
        RECT 139.800 111.800 140.200 112.200 ;
        RECT 3.000 105.800 3.400 106.200 ;
        RECT 5.400 106.800 5.800 107.200 ;
        RECT 16.600 108.800 17.000 109.200 ;
        RECT 6.200 105.800 6.600 106.200 ;
        RECT 8.600 105.800 9.000 106.200 ;
        RECT 2.200 103.800 2.600 104.200 ;
        RECT 11.800 103.800 12.200 104.200 ;
        RECT 8.600 101.800 9.000 102.200 ;
        RECT 12.600 101.800 13.000 102.200 ;
        RECT 15.000 104.800 15.400 105.200 ;
        RECT 14.200 101.800 14.600 102.200 ;
        RECT 27.000 108.800 27.400 109.200 ;
        RECT 21.400 105.800 21.800 106.200 ;
        RECT 19.000 104.800 19.400 105.200 ;
        RECT 24.600 105.800 25.000 106.200 ;
        RECT 25.400 105.800 25.800 106.200 ;
        RECT 27.800 106.800 28.200 107.200 ;
        RECT 36.600 108.800 37.000 109.200 ;
        RECT 39.800 108.800 40.200 109.200 ;
        RECT 18.200 101.800 18.600 102.200 ;
        RECT 21.400 102.800 21.800 103.200 ;
        RECT 37.400 106.800 37.800 107.200 ;
        RECT 38.200 105.800 38.600 106.200 ;
        RECT 40.600 106.800 41.000 107.200 ;
        RECT 61.400 108.800 61.800 109.200 ;
        RECT 60.600 106.800 61.000 107.200 ;
        RECT 48.600 105.800 49.000 106.200 ;
        RECT 59.000 105.800 59.400 106.200 ;
        RECT 66.200 108.800 66.600 109.200 ;
        RECT 64.600 106.800 65.000 107.200 ;
        RECT 80.600 108.800 81.000 109.200 ;
        RECT 55.000 103.800 55.400 104.200 ;
        RECT 65.400 104.800 65.800 105.200 ;
        RECT 71.000 105.800 71.400 106.200 ;
        RECT 74.200 106.800 74.600 107.200 ;
        RECT 75.000 105.800 75.400 106.200 ;
        RECT 78.200 107.800 78.600 108.200 ;
        RECT 79.800 107.800 80.200 108.200 ;
        RECT 77.400 104.800 77.800 105.200 ;
        RECT 81.400 106.800 81.800 107.200 ;
        RECT 87.000 108.800 87.400 109.200 ;
        RECT 82.200 105.800 82.600 106.200 ;
        RECT 83.800 104.800 84.200 105.200 ;
        RECT 89.400 108.800 89.800 109.200 ;
        RECT 92.600 108.800 93.000 109.200 ;
        RECT 88.600 106.800 89.000 107.200 ;
        RECT 91.800 106.800 92.200 107.200 ;
        RECT 107.000 106.500 107.400 106.900 ;
        RECT 102.200 105.800 102.600 106.200 ;
        RECT 87.000 101.800 87.400 102.200 ;
        RECT 111.800 106.300 112.200 106.700 ;
        RECT 115.000 105.800 115.400 106.200 ;
        RECT 107.800 104.400 108.200 104.800 ;
        RECT 110.200 103.800 110.600 104.200 ;
        RECT 108.600 103.100 109.000 103.500 ;
        RECT 107.000 102.100 107.400 102.500 ;
        RECT 107.800 102.100 108.200 102.500 ;
        RECT 110.200 103.100 110.600 103.500 ;
        RECT 111.800 103.100 112.200 103.500 ;
        RECT 112.600 102.100 113.000 102.500 ;
        RECT 113.400 102.100 113.800 102.500 ;
        RECT 114.200 102.100 114.600 102.500 ;
        RECT 127.800 106.500 128.200 106.900 ;
        RECT 119.000 101.800 119.400 102.200 ;
        RECT 132.600 106.300 133.000 106.700 ;
        RECT 124.600 105.800 125.000 106.200 ;
        RECT 127.000 105.800 127.400 106.200 ;
        RECT 128.600 104.400 129.000 104.800 ;
        RECT 131.000 103.800 131.400 104.200 ;
        RECT 129.400 103.100 129.800 103.500 ;
        RECT 127.800 102.100 128.200 102.500 ;
        RECT 128.600 102.100 129.000 102.500 ;
        RECT 131.000 103.100 131.400 103.500 ;
        RECT 132.600 103.100 133.000 103.500 ;
        RECT 133.400 102.100 133.800 102.500 ;
        RECT 134.200 102.100 134.600 102.500 ;
        RECT 135.000 102.100 135.400 102.500 ;
        RECT 140.600 103.800 141.000 104.200 ;
        RECT 147.800 105.800 148.200 106.200 ;
        RECT 2.200 98.800 2.600 99.200 ;
        RECT 1.400 96.800 1.800 97.200 ;
        RECT 3.000 95.800 3.400 96.200 ;
        RECT 3.800 93.800 4.200 94.200 ;
        RECT 7.000 98.800 7.400 99.200 ;
        RECT 6.200 96.800 6.600 97.200 ;
        RECT 7.800 95.800 8.200 96.200 ;
        RECT 7.000 94.800 7.400 95.200 ;
        RECT 4.600 91.800 5.000 92.200 ;
        RECT 8.600 93.800 9.000 94.200 ;
        RECT 16.600 98.800 17.000 99.200 ;
        RECT 15.800 96.800 16.200 97.200 ;
        RECT 11.000 94.800 11.400 95.200 ;
        RECT 17.400 95.800 17.800 96.200 ;
        RECT 16.600 94.800 17.000 95.200 ;
        RECT 22.200 94.800 22.600 95.200 ;
        RECT 29.400 98.800 29.800 99.200 ;
        RECT 32.600 98.800 33.000 99.200 ;
        RECT 28.600 96.800 29.000 97.200 ;
        RECT 31.800 96.800 32.200 97.200 ;
        RECT 30.200 95.800 30.600 96.200 ;
        RECT 29.400 94.800 29.800 95.200 ;
        RECT 33.400 95.800 33.800 96.200 ;
        RECT 39.000 96.800 39.400 97.200 ;
        RECT 46.200 98.800 46.600 99.200 ;
        RECT 51.000 98.800 51.400 99.200 ;
        RECT 40.600 96.800 41.000 97.200 ;
        RECT 37.400 95.800 37.800 96.200 ;
        RECT 32.600 94.800 33.000 95.200 ;
        RECT 25.400 91.800 25.800 92.200 ;
        RECT 43.800 96.800 44.200 97.200 ;
        RECT 47.000 96.800 47.400 97.200 ;
        RECT 51.800 96.800 52.200 97.200 ;
        RECT 55.000 96.800 55.400 97.200 ;
        RECT 59.000 98.800 59.400 99.200 ;
        RECT 62.200 98.800 62.600 99.200 ;
        RECT 42.200 95.800 42.600 96.200 ;
        RECT 45.400 95.800 45.800 96.200 ;
        RECT 50.200 95.800 50.600 96.200 ;
        RECT 53.400 95.800 53.800 96.200 ;
        RECT 59.800 96.800 60.200 97.200 ;
        RECT 41.400 93.800 41.800 94.200 ;
        RECT 61.400 95.800 61.800 96.200 ;
        RECT 65.400 98.800 65.800 99.200 ;
        RECT 69.400 98.800 69.800 99.200 ;
        RECT 70.200 96.800 70.600 97.200 ;
        RECT 60.600 94.800 61.000 95.200 ;
        RECT 68.600 95.800 69.000 96.200 ;
        RECT 83.000 98.800 83.400 99.200 ;
        RECT 58.200 92.800 58.600 93.200 ;
        RECT 67.800 93.800 68.200 94.200 ;
        RECT 91.000 98.800 91.400 99.200 ;
        RECT 79.800 94.800 80.200 95.200 ;
        RECT 95.800 96.800 96.200 97.200 ;
        RECT 106.200 98.800 106.600 99.200 ;
        RECT 77.400 93.800 77.800 94.200 ;
        RECT 83.800 93.800 84.200 94.200 ;
        RECT 91.000 94.800 91.400 95.200 ;
        RECT 97.400 95.800 97.800 96.200 ;
        RECT 102.200 95.800 102.600 96.200 ;
        RECT 96.600 94.800 97.000 95.200 ;
        RECT 99.000 94.800 99.400 95.200 ;
        RECT 103.800 94.800 104.200 95.200 ;
        RECT 88.600 93.800 89.000 94.200 ;
        RECT 91.800 93.800 92.200 94.200 ;
        RECT 94.200 92.800 94.600 93.200 ;
        RECT 120.600 98.800 121.000 99.200 ;
        RECT 109.400 92.800 109.800 93.200 ;
        RECT 111.800 92.800 112.200 93.200 ;
        RECT 115.800 94.800 116.200 95.200 ;
        RECT 114.200 93.800 114.600 94.200 ;
        RECT 121.400 92.800 121.800 93.200 ;
        RECT 132.600 97.500 133.000 97.900 ;
        RECT 131.000 96.800 131.400 97.200 ;
        RECT 133.400 96.200 133.800 96.600 ;
        RECT 127.800 94.100 128.200 94.500 ;
        RECT 132.600 94.300 133.000 94.700 ;
        RECT 130.200 93.800 130.600 94.200 ;
        RECT 139.900 94.800 140.300 95.200 ;
        RECT 127.800 92.100 128.200 92.500 ;
        RECT 128.600 92.100 129.000 92.500 ;
        RECT 129.400 92.100 129.800 92.500 ;
        RECT 131.000 92.100 131.400 92.500 ;
        RECT 132.600 92.100 133.000 92.500 ;
        RECT 133.400 92.100 133.800 92.500 ;
        RECT 134.200 92.100 134.600 92.500 ;
        RECT 135.000 92.100 135.400 92.500 ;
        RECT 146.200 94.800 146.600 95.200 ;
        RECT 143.800 92.800 144.200 93.200 ;
        RECT 148.600 92.800 149.000 93.200 ;
        RECT 149.400 91.800 149.800 92.200 ;
        RECT 3.800 88.800 4.200 89.200 ;
        RECT 1.400 86.800 1.800 87.200 ;
        RECT 7.800 88.800 8.200 89.200 ;
        RECT 8.600 85.800 9.000 86.200 ;
        RECT 14.200 88.800 14.600 89.200 ;
        RECT 11.800 86.800 12.200 87.200 ;
        RECT 22.200 88.800 22.600 89.200 ;
        RECT 12.600 85.800 13.000 86.200 ;
        RECT 15.000 85.800 15.400 86.200 ;
        RECT 3.000 81.800 3.400 82.200 ;
        RECT 24.600 86.800 25.000 87.200 ;
        RECT 15.800 83.800 16.200 84.200 ;
        RECT 43.800 88.800 44.200 89.200 ;
        RECT 63.800 88.800 64.200 89.200 ;
        RECT 30.200 85.800 30.600 86.200 ;
        RECT 35.800 85.800 36.200 86.200 ;
        RECT 39.000 86.800 39.400 87.200 ;
        RECT 39.800 85.800 40.200 86.200 ;
        RECT 32.600 83.800 33.000 84.200 ;
        RECT 43.000 84.800 43.400 85.200 ;
        RECT 47.800 85.800 48.200 86.200 ;
        RECT 51.800 84.800 52.200 85.200 ;
        RECT 55.000 84.800 55.400 85.200 ;
        RECT 67.000 88.800 67.400 89.200 ;
        RECT 70.200 86.800 70.600 87.200 ;
        RECT 71.800 86.800 72.200 87.200 ;
        RECT 69.400 85.800 69.800 86.200 ;
        RECT 72.600 84.800 73.000 85.200 ;
        RECT 79.000 88.800 79.400 89.200 ;
        RECT 83.800 88.800 84.200 89.200 ;
        RECT 84.600 88.800 85.000 89.200 ;
        RECT 79.000 87.400 79.400 87.800 ;
        RECT 80.600 86.800 81.000 87.200 ;
        RECT 84.600 81.800 85.000 82.200 ;
        RECT 87.000 87.800 87.400 88.200 ;
        RECT 92.600 88.800 93.000 89.200 ;
        RECT 91.800 86.800 92.200 87.200 ;
        RECT 93.400 86.800 93.800 87.200 ;
        RECT 91.000 84.800 91.400 85.200 ;
        RECT 96.600 85.800 97.000 86.200 ;
        RECT 103.800 87.400 104.200 87.800 ;
        RECT 105.400 86.800 105.800 87.200 ;
        RECT 112.600 88.800 113.000 89.200 ;
        RECT 111.800 86.800 112.200 87.200 ;
        RECT 109.400 81.800 109.800 82.200 ;
        RECT 116.600 85.800 117.000 86.200 ;
        RECT 124.600 88.800 125.000 89.200 ;
        RECT 123.000 86.800 123.400 87.200 ;
        RECT 123.800 86.800 124.200 87.200 ;
        RECT 127.800 86.800 128.200 87.200 ;
        RECT 134.200 87.400 134.600 87.800 ;
        RECT 131.000 86.800 131.400 87.200 ;
        RECT 130.200 85.800 130.600 86.200 ;
        RECT 128.600 84.800 129.000 85.200 ;
        RECT 139.800 88.800 140.200 89.200 ;
        RECT 141.400 88.800 141.800 89.200 ;
        RECT 137.400 86.800 137.800 87.200 ;
        RECT 139.000 86.800 139.400 87.200 ;
        RECT 131.800 84.800 132.200 85.200 ;
        RECT 135.800 85.800 136.200 86.200 ;
        RECT 148.600 84.800 149.000 85.200 ;
        RECT 149.400 81.800 149.800 82.200 ;
        RECT 2.200 78.800 2.600 79.200 ;
        RECT 1.400 76.800 1.800 77.200 ;
        RECT 7.800 76.800 8.200 77.200 ;
        RECT 3.000 75.800 3.400 76.200 ;
        RECT 2.200 74.800 2.600 75.200 ;
        RECT 5.400 74.800 5.800 75.200 ;
        RECT 9.400 75.800 9.800 76.200 ;
        RECT 15.800 78.800 16.200 79.200 ;
        RECT 15.000 76.800 15.400 77.200 ;
        RECT 13.400 75.800 13.800 76.200 ;
        RECT 8.600 74.800 9.000 75.200 ;
        RECT 4.600 73.800 5.000 74.200 ;
        RECT 6.200 73.800 6.600 74.200 ;
        RECT 19.800 74.800 20.200 75.200 ;
        RECT 23.000 74.800 23.400 75.200 ;
        RECT 18.200 73.800 18.600 74.200 ;
        RECT 17.400 72.800 17.800 73.200 ;
        RECT 27.000 73.800 27.400 74.200 ;
        RECT 26.200 72.800 26.600 73.200 ;
        RECT 27.800 72.800 28.200 73.200 ;
        RECT 33.400 74.800 33.800 75.200 ;
        RECT 31.800 73.800 32.200 74.200 ;
        RECT 42.200 76.800 42.600 77.200 ;
        RECT 50.200 78.800 50.600 79.200 ;
        RECT 51.000 76.800 51.400 77.200 ;
        RECT 52.600 77.800 53.000 78.200 ;
        RECT 55.000 78.800 55.400 79.200 ;
        RECT 49.400 75.800 49.800 76.200 ;
        RECT 45.400 72.800 45.800 73.200 ;
        RECT 55.800 76.800 56.200 77.200 ;
        RECT 59.000 76.800 59.400 77.200 ;
        RECT 64.600 78.800 65.000 79.200 ;
        RECT 77.400 78.800 77.800 79.200 ;
        RECT 76.600 76.800 77.000 77.200 ;
        RECT 72.600 74.800 73.000 75.200 ;
        RECT 53.400 72.800 53.800 73.200 ;
        RECT 66.200 73.800 66.600 74.200 ;
        RECT 62.200 72.800 62.600 73.200 ;
        RECT 69.400 72.800 69.800 73.200 ;
        RECT 75.000 73.800 75.400 74.200 ;
        RECT 76.600 73.800 77.000 74.200 ;
        RECT 82.200 78.800 82.600 79.200 ;
        RECT 87.800 78.800 88.200 79.200 ;
        RECT 81.400 73.800 81.800 74.200 ;
        RECT 90.200 74.800 90.600 75.200 ;
        RECT 87.000 73.800 87.400 74.200 ;
        RECT 78.200 71.800 78.600 72.200 ;
        RECT 79.800 71.800 80.200 72.200 ;
        RECT 92.600 73.800 93.000 74.200 ;
        RECT 88.600 72.800 89.000 73.200 ;
        RECT 103.800 78.800 104.200 79.200 ;
        RECT 103.000 73.800 103.400 74.200 ;
        RECT 91.800 71.800 92.200 72.200 ;
        RECT 111.000 78.800 111.400 79.200 ;
        RECT 119.000 78.800 119.400 79.200 ;
        RECT 104.600 72.800 105.000 73.200 ;
        RECT 106.200 71.800 106.600 72.200 ;
        RECT 121.400 75.800 121.800 76.200 ;
        RECT 119.000 74.800 119.400 75.200 ;
        RECT 128.600 77.800 129.000 78.200 ;
        RECT 110.200 71.800 110.600 72.200 ;
        RECT 116.600 72.800 117.000 73.200 ;
        RECT 122.200 73.800 122.600 74.200 ;
        RECT 132.600 75.800 133.000 76.200 ;
        RECT 141.400 78.800 141.800 79.200 ;
        RECT 131.800 73.800 132.200 74.200 ;
        RECT 123.800 71.800 124.200 72.200 ;
        RECT 134.200 74.800 134.600 75.200 ;
        RECT 137.400 74.800 137.800 75.200 ;
        RECT 146.200 78.800 146.600 79.200 ;
        RECT 141.400 74.800 141.800 75.200 ;
        RECT 142.200 73.800 142.600 74.200 ;
        RECT 143.000 72.800 143.400 73.200 ;
        RECT 150.200 75.800 150.600 76.200 ;
        RECT 146.200 71.800 146.600 72.200 ;
        RECT 1.400 66.800 1.800 67.200 ;
        RECT 7.800 66.800 8.200 67.200 ;
        RECT 8.600 65.800 9.000 66.200 ;
        RECT 14.200 65.800 14.600 66.200 ;
        RECT 31.800 68.800 32.200 69.200 ;
        RECT 39.000 68.800 39.400 69.200 ;
        RECT 44.600 68.800 45.000 69.200 ;
        RECT 45.400 68.800 45.800 69.200 ;
        RECT 52.600 68.800 53.000 69.200 ;
        RECT 64.600 68.800 65.000 69.200 ;
        RECT 21.400 66.800 21.800 67.200 ;
        RECT 22.200 65.800 22.600 66.200 ;
        RECT 16.600 63.800 17.000 64.200 ;
        RECT 42.200 66.800 42.600 67.200 ;
        RECT 50.200 66.800 50.600 67.200 ;
        RECT 43.000 65.800 43.400 66.200 ;
        RECT 45.400 64.800 45.800 65.200 ;
        RECT 51.000 65.800 51.400 66.200 ;
        RECT 52.600 64.800 53.000 65.200 ;
        RECT 59.800 66.800 60.200 67.200 ;
        RECT 63.000 65.800 63.400 66.200 ;
        RECT 68.600 68.800 69.000 69.200 ;
        RECT 65.400 66.800 65.800 67.200 ;
        RECT 73.400 68.800 73.800 69.200 ;
        RECT 84.600 68.800 85.000 69.200 ;
        RECT 87.000 68.800 87.400 69.200 ;
        RECT 77.400 64.800 77.800 65.200 ;
        RECT 80.600 61.800 81.000 62.200 ;
        RECT 84.600 64.800 85.000 65.200 ;
        RECT 87.000 64.800 87.400 65.200 ;
        RECT 91.800 65.800 92.200 66.200 ;
        RECT 94.200 64.800 94.600 65.200 ;
        RECT 96.600 65.800 97.000 66.200 ;
        RECT 104.600 65.800 105.000 66.200 ;
        RECT 103.800 64.800 104.200 65.200 ;
        RECT 122.200 67.800 122.600 68.200 ;
        RECT 117.400 66.800 117.800 67.200 ;
        RECT 121.400 66.800 121.800 67.200 ;
        RECT 106.200 64.800 106.600 65.200 ;
        RECT 108.600 61.800 109.000 62.200 ;
        RECT 118.200 64.800 118.600 65.200 ;
        RECT 120.600 65.800 121.000 66.200 ;
        RECT 123.000 64.800 123.400 65.200 ;
        RECT 130.200 68.800 130.600 69.200 ;
        RECT 131.800 67.800 132.200 68.200 ;
        RECT 143.000 68.800 143.400 69.200 ;
        RECT 143.800 68.800 144.200 69.200 ;
        RECT 130.200 64.800 130.600 65.200 ;
        RECT 133.400 66.800 133.800 67.200 ;
        RECT 139.000 66.800 139.400 67.200 ;
        RECT 135.800 65.800 136.200 66.200 ;
        RECT 136.600 65.800 137.000 66.200 ;
        RECT 139.800 65.800 140.200 66.200 ;
        RECT 137.400 64.800 137.800 65.200 ;
        RECT 145.400 66.800 145.800 67.200 ;
        RECT 148.600 66.800 149.000 67.200 ;
        RECT 149.400 65.800 149.800 66.200 ;
        RECT 3.800 56.800 4.200 57.200 ;
        RECT 0.600 52.800 1.000 53.200 ;
        RECT 13.400 58.800 13.800 59.200 ;
        RECT 19.000 58.800 19.400 59.200 ;
        RECT 21.400 58.800 21.800 59.200 ;
        RECT 19.800 56.800 20.200 57.200 ;
        RECT 22.200 56.800 22.600 57.200 ;
        RECT 25.400 56.800 25.800 57.200 ;
        RECT 13.400 54.800 13.800 55.200 ;
        RECT 18.200 55.800 18.600 56.200 ;
        RECT 7.000 53.800 7.400 54.200 ;
        RECT 7.800 52.800 8.200 53.200 ;
        RECT 11.000 53.800 11.400 54.200 ;
        RECT 14.200 53.800 14.600 54.200 ;
        RECT 23.800 55.800 24.200 56.200 ;
        RECT 23.000 54.800 23.400 55.200 ;
        RECT 27.000 55.800 27.400 56.200 ;
        RECT 35.000 58.800 35.400 59.200 ;
        RECT 32.600 56.800 33.000 57.200 ;
        RECT 35.800 56.800 36.200 57.200 ;
        RECT 31.000 55.800 31.400 56.200 ;
        RECT 34.200 55.800 34.600 56.200 ;
        RECT 26.200 54.800 26.600 55.200 ;
        RECT 8.600 51.800 9.000 52.200 ;
        RECT 16.600 51.800 17.000 52.200 ;
        RECT 38.200 54.800 38.600 55.200 ;
        RECT 39.800 54.800 40.200 55.200 ;
        RECT 57.400 58.800 57.800 59.200 ;
        RECT 61.400 58.800 61.800 59.200 ;
        RECT 28.600 51.800 29.000 52.200 ;
        RECT 41.400 53.800 41.800 54.200 ;
        RECT 46.200 52.800 46.600 53.200 ;
        RECT 51.000 53.800 51.400 54.200 ;
        RECT 55.000 52.800 55.400 53.200 ;
        RECT 60.600 53.800 61.000 54.200 ;
        RECT 63.800 58.800 64.200 59.200 ;
        RECT 63.000 53.800 63.400 54.200 ;
        RECT 63.800 51.800 64.200 52.200 ;
        RECT 67.000 52.800 67.400 53.200 ;
        RECT 69.400 52.800 69.800 53.200 ;
        RECT 67.800 51.800 68.200 52.200 ;
        RECT 75.000 52.800 75.400 53.200 ;
        RECT 79.000 56.800 79.400 57.200 ;
        RECT 79.800 53.800 80.200 54.200 ;
        RECT 86.200 54.800 86.600 55.200 ;
        RECT 75.800 51.800 76.200 52.200 ;
        RECT 83.800 51.800 84.200 52.200 ;
        RECT 91.000 54.800 91.400 55.200 ;
        RECT 94.200 54.800 94.600 55.200 ;
        RECT 101.400 54.800 101.800 55.200 ;
        RECT 89.400 51.800 89.800 52.200 ;
        RECT 92.600 51.800 93.000 52.200 ;
        RECT 105.400 53.800 105.800 54.200 ;
        RECT 103.800 52.800 104.200 53.200 ;
        RECT 105.400 52.800 105.800 53.200 ;
        RECT 111.800 54.800 112.200 55.200 ;
        RECT 108.600 51.800 109.000 52.200 ;
        RECT 116.600 54.800 117.000 55.200 ;
        RECT 119.000 53.800 119.400 54.200 ;
        RECT 130.200 56.800 130.600 57.200 ;
        RECT 135.800 58.800 136.200 59.200 ;
        RECT 135.000 56.800 135.400 57.200 ;
        RECT 115.000 51.800 115.400 52.200 ;
        RECT 127.800 54.800 128.200 55.200 ;
        RECT 133.400 55.800 133.800 56.200 ;
        RECT 123.000 52.800 123.400 53.200 ;
        RECT 125.400 52.800 125.800 53.200 ;
        RECT 136.600 53.800 137.000 54.200 ;
        RECT 144.600 54.800 145.000 55.200 ;
        RECT 141.400 53.800 141.800 54.200 ;
        RECT 137.400 51.800 137.800 52.200 ;
        RECT 142.200 52.800 142.600 53.200 ;
        RECT 147.800 52.800 148.200 53.200 ;
        RECT 148.600 52.800 149.000 53.200 ;
        RECT 149.400 51.800 149.800 52.200 ;
        RECT 2.200 46.600 2.600 47.000 ;
        RECT 3.000 46.800 3.400 47.200 ;
        RECT 0.600 41.800 1.000 42.200 ;
        RECT 7.800 45.800 8.200 46.200 ;
        RECT 5.400 44.800 5.800 45.200 ;
        RECT 7.800 43.800 8.200 44.200 ;
        RECT 11.000 44.800 11.400 45.200 ;
        RECT 16.600 45.800 17.000 46.200 ;
        RECT 15.800 44.800 16.200 45.200 ;
        RECT 25.400 48.800 25.800 49.200 ;
        RECT 22.200 47.400 22.600 47.800 ;
        RECT 37.400 48.800 37.800 49.200 ;
        RECT 23.800 46.800 24.200 47.200 ;
        RECT 31.800 46.800 32.200 47.200 ;
        RECT 34.200 46.800 34.600 47.200 ;
        RECT 35.800 46.800 36.200 47.200 ;
        RECT 57.400 48.800 57.800 49.200 ;
        RECT 27.000 45.800 27.400 46.200 ;
        RECT 21.400 41.800 21.800 42.200 ;
        RECT 35.000 45.800 35.400 46.200 ;
        RECT 36.600 44.800 37.000 45.200 ;
        RECT 40.600 45.800 41.000 46.200 ;
        RECT 45.400 45.800 45.800 46.200 ;
        RECT 52.600 45.800 53.000 46.200 ;
        RECT 64.600 48.800 65.000 49.200 ;
        RECT 70.200 46.800 70.600 47.200 ;
        RECT 62.200 41.800 62.600 42.200 ;
        RECT 68.600 41.800 69.000 42.200 ;
        RECT 71.000 41.800 71.400 42.200 ;
        RECT 104.600 48.800 105.000 49.200 ;
        RECT 82.200 46.800 82.600 47.200 ;
        RECT 87.800 46.800 88.200 47.200 ;
        RECT 93.400 46.800 93.800 47.200 ;
        RECT 78.200 45.800 78.600 46.200 ;
        RECT 84.600 45.800 85.000 46.200 ;
        RECT 85.400 45.800 85.800 46.200 ;
        RECT 73.400 41.800 73.800 42.200 ;
        RECT 76.600 41.800 77.000 42.200 ;
        RECT 83.000 44.800 83.400 45.200 ;
        RECT 86.200 44.800 86.600 45.200 ;
        RECT 93.400 44.800 93.800 45.200 ;
        RECT 100.600 46.800 101.000 47.200 ;
        RECT 99.800 45.800 100.200 46.200 ;
        RECT 99.000 44.800 99.400 45.200 ;
        RECT 102.200 41.800 102.600 42.200 ;
        RECT 110.200 44.800 110.600 45.200 ;
        RECT 120.600 46.800 121.000 47.200 ;
        RECT 115.000 45.800 115.400 46.200 ;
        RECT 111.000 41.800 111.400 42.200 ;
        RECT 117.400 44.800 117.800 45.200 ;
        RECT 124.600 46.800 125.000 47.200 ;
        RECT 120.600 44.800 121.000 45.200 ;
        RECT 121.400 44.800 121.800 45.200 ;
        RECT 127.000 45.800 127.400 46.200 ;
        RECT 131.800 44.800 132.200 45.200 ;
        RECT 131.000 41.800 131.400 42.200 ;
        RECT 138.200 48.800 138.600 49.200 ;
        RECT 136.600 45.800 137.000 46.200 ;
        RECT 133.400 41.800 133.800 42.200 ;
        RECT 136.600 43.800 137.000 44.200 ;
        RECT 141.400 48.800 141.800 49.200 ;
        RECT 139.800 46.800 140.200 47.200 ;
        RECT 140.600 46.800 141.000 47.200 ;
        RECT 143.000 44.800 143.400 45.200 ;
        RECT 150.200 45.800 150.600 46.200 ;
        RECT 2.200 38.800 2.600 39.200 ;
        RECT 7.800 38.800 8.200 39.200 ;
        RECT 8.600 36.800 9.000 37.200 ;
        RECT 14.200 38.800 14.600 39.200 ;
        RECT 2.200 34.800 2.600 35.200 ;
        RECT 7.000 35.800 7.400 36.200 ;
        RECT 15.000 36.800 15.400 37.200 ;
        RECT 3.000 33.800 3.400 34.200 ;
        RECT 11.000 34.800 11.400 35.200 ;
        RECT 13.400 35.800 13.800 36.200 ;
        RECT 20.600 38.800 21.000 39.200 ;
        RECT 21.400 36.800 21.800 37.200 ;
        RECT 19.800 35.800 20.200 36.200 ;
        RECT 23.900 35.900 24.300 36.300 ;
        RECT 24.500 34.900 24.900 35.300 ;
        RECT 23.900 33.100 24.300 33.500 ;
        RECT 27.800 33.800 28.200 34.200 ;
        RECT 31.000 38.800 31.400 39.200 ;
        RECT 34.200 38.800 34.600 39.200 ;
        RECT 36.600 38.800 37.000 39.200 ;
        RECT 31.800 32.800 32.200 33.200 ;
        RECT 39.800 38.800 40.200 39.200 ;
        RECT 42.200 36.800 42.600 37.200 ;
        RECT 37.400 33.800 37.800 34.200 ;
        RECT 36.600 32.800 37.000 33.200 ;
        RECT 57.400 37.800 57.800 38.200 ;
        RECT 61.400 38.800 61.800 39.200 ;
        RECT 47.000 33.800 47.400 34.200 ;
        RECT 55.000 33.800 55.400 34.200 ;
        RECT 59.000 34.800 59.400 35.200 ;
        RECT 59.800 34.800 60.200 35.200 ;
        RECT 74.200 38.800 74.600 39.200 ;
        RECT 77.400 36.800 77.800 37.200 ;
        RECT 85.400 38.800 85.800 39.200 ;
        RECT 68.600 34.800 69.000 35.200 ;
        RECT 69.400 34.800 69.800 35.200 ;
        RECT 70.200 34.800 70.600 35.200 ;
        RECT 66.200 32.800 66.600 33.200 ;
        RECT 75.800 34.800 76.200 35.200 ;
        RECT 79.800 34.800 80.200 35.200 ;
        RECT 82.200 34.800 82.600 35.200 ;
        RECT 80.600 33.800 81.000 34.200 ;
        RECT 78.200 31.800 78.600 32.200 ;
        RECT 83.800 32.800 84.200 33.200 ;
        RECT 88.600 36.800 89.000 37.200 ;
        RECT 86.200 33.800 86.600 34.200 ;
        RECT 87.000 32.800 87.400 33.200 ;
        RECT 95.800 34.800 96.200 35.200 ;
        RECT 105.400 37.800 105.800 38.200 ;
        RECT 94.200 32.800 94.600 33.200 ;
        RECT 101.400 34.800 101.800 35.200 ;
        RECT 102.200 33.800 102.600 34.200 ;
        RECT 104.600 33.800 105.000 34.200 ;
        RECT 97.400 31.800 97.800 32.200 ;
        RECT 99.000 31.800 99.400 32.200 ;
        RECT 108.600 37.800 109.000 38.200 ;
        RECT 109.400 34.800 109.800 35.200 ;
        RECT 106.200 33.800 106.600 34.200 ;
        RECT 109.400 33.800 109.800 34.200 ;
        RECT 111.800 32.800 112.200 33.200 ;
        RECT 119.000 33.800 119.400 34.200 ;
        RECT 133.400 38.800 133.800 39.200 ;
        RECT 115.000 31.800 115.400 32.200 ;
        RECT 118.200 31.800 118.600 32.200 ;
        RECT 121.400 32.800 121.800 33.200 ;
        RECT 131.800 33.800 132.200 34.200 ;
        RECT 132.600 32.800 133.000 33.200 ;
        RECT 136.600 38.800 137.000 39.200 ;
        RECT 135.800 36.800 136.200 37.200 ;
        RECT 137.400 35.800 137.800 36.200 ;
        RECT 136.600 34.800 137.000 35.200 ;
        RECT 134.200 33.800 134.600 34.200 ;
        RECT 139.800 33.800 140.200 34.200 ;
        RECT 141.400 32.800 141.800 33.200 ;
        RECT 146.200 31.800 146.600 32.200 ;
        RECT 3.800 27.400 4.200 27.800 ;
        RECT 7.000 28.800 7.400 29.200 ;
        RECT 11.000 28.800 11.400 29.200 ;
        RECT 5.400 26.800 5.800 27.200 ;
        RECT 10.200 26.800 10.600 27.200 ;
        RECT 7.800 25.800 8.200 26.200 ;
        RECT 15.000 28.800 15.400 29.200 ;
        RECT 14.200 26.800 14.600 27.200 ;
        RECT 3.800 23.800 4.200 24.200 ;
        RECT 8.600 23.800 9.000 24.200 ;
        RECT 15.800 26.800 16.200 27.200 ;
        RECT 16.600 25.800 17.000 26.200 ;
        RECT 22.200 26.800 22.600 27.200 ;
        RECT 51.800 28.800 52.200 29.200 ;
        RECT 24.600 21.800 25.000 22.200 ;
        RECT 27.800 21.800 28.200 22.200 ;
        RECT 34.200 24.800 34.600 25.200 ;
        RECT 39.800 21.800 40.200 22.200 ;
        RECT 43.800 21.800 44.200 22.200 ;
        RECT 63.000 28.800 63.400 29.200 ;
        RECT 58.200 25.800 58.600 26.200 ;
        RECT 55.000 24.800 55.400 25.200 ;
        RECT 59.000 24.800 59.400 25.200 ;
        RECT 64.600 27.800 65.000 28.200 ;
        RECT 71.000 28.800 71.400 29.200 ;
        RECT 74.200 28.800 74.600 29.200 ;
        RECT 63.800 24.800 64.200 25.200 ;
        RECT 79.800 28.800 80.200 29.200 ;
        RECT 71.000 24.800 71.400 25.200 ;
        RECT 76.600 25.800 77.000 26.200 ;
        RECT 77.400 21.800 77.800 22.200 ;
        RECT 82.200 28.800 82.600 29.200 ;
        RECT 81.400 26.800 81.800 27.200 ;
        RECT 86.200 28.800 86.600 29.200 ;
        RECT 87.800 26.800 88.200 27.200 ;
        RECT 95.800 28.800 96.200 29.200 ;
        RECT 86.200 24.800 86.600 25.200 ;
        RECT 89.400 25.800 89.800 26.200 ;
        RECT 95.000 26.800 95.400 27.200 ;
        RECT 91.800 25.800 92.200 26.200 ;
        RECT 103.800 28.800 104.200 29.200 ;
        RECT 99.800 26.800 100.200 27.200 ;
        RECT 101.400 26.800 101.800 27.200 ;
        RECT 99.000 24.800 99.400 25.200 ;
        RECT 111.000 28.800 111.400 29.200 ;
        RECT 117.400 28.800 117.800 29.200 ;
        RECT 110.200 26.800 110.600 27.200 ;
        RECT 113.400 26.800 113.800 27.200 ;
        RECT 116.600 26.800 117.000 27.200 ;
        RECT 107.800 24.800 108.200 25.200 ;
        RECT 104.600 21.800 105.000 22.200 ;
        RECT 138.200 28.800 138.600 29.200 ;
        RECT 140.600 28.800 141.000 29.200 ;
        RECT 130.200 26.800 130.600 27.200 ;
        RECT 137.400 26.800 137.800 27.200 ;
        RECT 131.000 25.800 131.400 26.200 ;
        RECT 135.800 24.800 136.200 25.200 ;
        RECT 150.200 28.800 150.600 29.200 ;
        RECT 146.200 25.800 146.600 26.200 ;
        RECT 2.200 18.800 2.600 19.200 ;
        RECT 8.600 18.800 9.000 19.200 ;
        RECT 1.400 16.800 1.800 17.200 ;
        RECT 4.600 16.800 5.000 17.200 ;
        RECT 3.000 15.800 3.400 16.200 ;
        RECT 6.200 15.800 6.600 16.200 ;
        RECT 15.000 17.800 15.400 18.200 ;
        RECT 2.200 14.800 2.600 15.200 ;
        RECT 5.400 14.800 5.800 15.200 ;
        RECT 19.800 18.800 20.200 19.200 ;
        RECT 20.600 16.800 21.000 17.200 ;
        RECT 24.600 16.800 25.000 17.200 ;
        RECT 9.400 13.800 9.800 14.200 ;
        RECT 17.400 14.800 17.800 15.200 ;
        RECT 18.200 14.800 18.600 15.200 ;
        RECT 23.000 15.800 23.400 16.200 ;
        RECT 21.400 14.800 21.800 15.200 ;
        RECT 15.800 13.800 16.200 14.200 ;
        RECT 29.400 13.800 29.800 14.200 ;
        RECT 34.200 16.800 34.600 17.200 ;
        RECT 35.800 16.800 36.200 17.200 ;
        RECT 37.400 15.800 37.800 16.200 ;
        RECT 36.600 14.800 37.000 15.200 ;
        RECT 27.000 11.800 27.400 12.200 ;
        RECT 59.800 18.800 60.200 19.200 ;
        RECT 41.400 12.800 41.800 13.200 ;
        RECT 39.000 11.800 39.400 12.200 ;
        RECT 45.400 13.800 45.800 14.200 ;
        RECT 47.000 11.800 47.400 12.200 ;
        RECT 61.400 14.800 61.800 15.200 ;
        RECT 63.800 14.800 64.200 15.200 ;
        RECT 52.600 11.800 53.000 12.200 ;
        RECT 67.000 14.800 67.400 15.200 ;
        RECT 65.400 12.800 65.800 13.200 ;
        RECT 79.800 18.800 80.200 19.200 ;
        RECT 81.300 15.900 81.700 16.300 ;
        RECT 75.000 14.800 75.400 15.200 ;
        RECT 70.200 13.800 70.600 14.200 ;
        RECT 68.600 11.800 69.000 12.200 ;
        RECT 76.600 12.800 77.000 13.200 ;
        RECT 86.200 14.800 86.600 15.200 ;
        RECT 81.300 13.100 81.700 13.500 ;
        RECT 87.800 14.800 88.200 15.200 ;
        RECT 93.400 18.800 93.800 19.200 ;
        RECT 85.400 13.800 85.800 14.200 ;
        RECT 88.600 13.800 89.000 14.200 ;
        RECT 89.400 13.800 89.800 14.200 ;
        RECT 90.200 13.800 90.600 14.200 ;
        RECT 86.200 11.800 86.600 12.200 ;
        RECT 107.000 16.800 107.400 17.200 ;
        RECT 115.800 16.800 116.200 17.200 ;
        RECT 95.800 14.800 96.200 15.200 ;
        RECT 104.600 14.800 105.000 15.200 ;
        RECT 105.400 14.800 105.800 15.200 ;
        RECT 111.800 14.800 112.200 15.200 ;
        RECT 113.400 14.800 113.800 15.200 ;
        RECT 123.000 18.800 123.400 19.200 ;
        RECT 102.200 12.800 102.600 13.200 ;
        RECT 109.400 13.800 109.800 14.200 ;
        RECT 114.200 13.800 114.600 14.200 ;
        RECT 111.800 11.800 112.200 12.200 ;
        RECT 116.600 12.800 117.000 13.200 ;
        RECT 120.600 13.800 121.000 14.200 ;
        RECT 126.200 18.800 126.600 19.200 ;
        RECT 127.800 16.800 128.200 17.200 ;
        RECT 127.000 14.800 127.400 15.200 ;
        RECT 124.600 12.800 125.000 13.200 ;
        RECT 133.400 16.800 133.800 17.200 ;
        RECT 131.800 15.800 132.200 16.200 ;
        RECT 146.200 18.800 146.600 19.200 ;
        RECT 133.400 14.800 133.800 15.200 ;
        RECT 138.200 14.800 138.600 15.200 ;
        RECT 135.000 13.800 135.400 14.200 ;
        RECT 139.800 14.800 140.200 15.200 ;
        RECT 131.000 12.800 131.400 13.200 ;
        RECT 135.000 12.800 135.400 13.200 ;
        RECT 140.600 13.800 141.000 14.200 ;
        RECT 143.000 12.800 143.400 13.200 ;
        RECT 3.000 8.800 3.400 9.200 ;
        RECT 2.200 7.400 2.600 7.800 ;
        RECT 5.400 6.800 5.800 7.200 ;
        RECT 11.800 6.800 12.200 7.200 ;
        RECT 16.600 7.800 17.000 8.200 ;
        RECT 20.600 8.800 21.000 9.200 ;
        RECT 17.400 6.800 17.800 7.200 ;
        RECT 24.600 8.800 25.000 9.200 ;
        RECT 21.400 7.400 21.800 7.800 ;
        RECT 23.000 6.800 23.400 7.200 ;
        RECT 15.000 5.800 15.400 6.200 ;
        RECT 25.400 8.800 25.800 9.200 ;
        RECT 33.400 6.800 33.800 7.200 ;
        RECT 49.400 8.800 49.800 9.200 ;
        RECT 44.600 6.800 45.000 7.200 ;
        RECT 47.000 6.800 47.400 7.200 ;
        RECT 47.800 5.800 48.200 6.200 ;
        RECT 56.600 6.800 57.000 7.200 ;
        RECT 61.400 8.800 61.800 9.200 ;
        RECT 64.600 8.800 65.000 9.200 ;
        RECT 69.400 7.800 69.800 8.200 ;
        RECT 71.800 8.800 72.200 9.200 ;
        RECT 78.200 4.800 78.600 5.200 ;
        RECT 81.400 4.800 81.800 5.200 ;
        RECT 95.800 8.800 96.200 9.200 ;
        RECT 92.600 6.800 93.000 7.200 ;
        RECT 95.000 6.800 95.400 7.200 ;
        RECT 102.200 6.800 102.600 7.200 ;
        RECT 84.600 5.800 85.000 6.200 ;
        RECT 86.200 5.800 86.600 6.200 ;
        RECT 99.000 5.800 99.400 6.200 ;
        RECT 107.800 4.800 108.200 5.200 ;
        RECT 119.000 8.800 119.400 9.200 ;
        RECT 115.800 6.800 116.200 7.200 ;
        RECT 110.200 5.800 110.600 6.200 ;
        RECT 127.800 7.800 128.200 8.200 ;
        RECT 132.600 6.800 133.000 7.200 ;
        RECT 137.400 6.800 137.800 7.200 ;
        RECT 130.200 5.800 130.600 6.200 ;
        RECT 132.600 5.800 133.000 6.200 ;
        RECT 131.800 4.800 132.200 5.200 ;
        RECT 141.400 8.800 141.800 9.200 ;
        RECT 144.600 8.800 145.000 9.200 ;
        RECT 143.800 6.800 144.200 7.200 ;
        RECT 147.800 6.800 148.200 7.200 ;
        RECT 149.400 4.800 149.800 5.200 ;
      LAYER metal2 ;
        RECT 10.200 128.800 10.600 129.200 ;
        RECT 46.200 129.100 46.600 129.200 ;
        RECT 47.000 129.100 47.400 129.200 ;
        RECT 46.200 128.800 47.400 129.100 ;
        RECT 6.200 127.800 6.600 128.200 ;
        RECT 7.000 127.800 7.400 128.200 ;
        RECT 0.600 126.800 1.000 127.200 ;
        RECT 1.400 126.800 1.800 127.200 ;
        RECT 3.800 127.100 4.200 127.200 ;
        RECT 4.600 127.100 5.000 127.200 ;
        RECT 3.800 126.800 5.000 127.100 ;
        RECT 0.600 126.200 0.900 126.800 ;
        RECT 0.600 125.800 1.000 126.200 ;
        RECT 1.400 124.200 1.700 126.800 ;
        RECT 2.200 125.800 2.600 126.200 ;
        RECT 3.800 125.800 4.200 126.200 ;
        RECT 2.200 124.200 2.500 125.800 ;
        RECT 3.000 124.800 3.400 125.200 ;
        RECT 1.400 123.800 1.800 124.200 ;
        RECT 2.200 123.800 2.600 124.200 ;
        RECT 1.400 123.100 1.700 123.800 ;
        RECT 1.400 122.800 2.500 123.100 ;
        RECT 2.200 119.200 2.500 122.800 ;
        RECT 3.000 121.200 3.300 124.800 ;
        RECT 3.800 124.200 4.100 125.800 ;
        RECT 3.800 123.800 4.200 124.200 ;
        RECT 6.200 121.200 6.500 127.800 ;
        RECT 7.000 127.200 7.300 127.800 ;
        RECT 7.000 126.800 7.400 127.200 ;
        RECT 8.600 126.800 9.000 127.200 ;
        RECT 9.400 126.800 9.800 127.200 ;
        RECT 8.600 125.200 8.900 126.800 ;
        RECT 9.400 126.200 9.700 126.800 ;
        RECT 9.400 125.800 9.800 126.200 ;
        RECT 10.200 125.200 10.500 128.800 ;
        RECT 13.400 127.800 13.800 128.200 ;
        RECT 23.800 127.800 24.200 128.200 ;
        RECT 27.000 127.800 27.400 128.200 ;
        RECT 27.800 127.800 28.200 128.200 ;
        RECT 31.800 127.800 32.200 128.200 ;
        RECT 40.600 127.800 41.000 128.200 ;
        RECT 47.800 127.800 48.200 128.200 ;
        RECT 56.600 128.100 57.000 128.200 ;
        RECT 57.400 128.100 57.800 128.200 ;
        RECT 56.600 127.800 57.800 128.100 ;
        RECT 61.400 127.800 61.800 128.200 ;
        RECT 62.200 127.800 62.600 128.200 ;
        RECT 65.400 128.100 65.800 128.200 ;
        RECT 66.200 128.100 66.600 128.200 ;
        RECT 65.400 127.800 66.600 128.100 ;
        RECT 71.800 127.800 72.200 128.200 ;
        RECT 13.400 127.200 13.700 127.800 ;
        RECT 13.400 126.800 13.800 127.200 ;
        RECT 14.200 126.800 14.600 127.200 ;
        RECT 15.000 127.100 15.400 127.200 ;
        RECT 15.800 127.100 16.200 127.200 ;
        RECT 15.000 126.800 16.200 127.100 ;
        RECT 18.200 126.800 18.600 127.200 ;
        RECT 19.800 127.100 20.200 127.200 ;
        RECT 20.600 127.100 21.000 127.200 ;
        RECT 19.800 126.800 21.000 127.100 ;
        RECT 14.200 126.200 14.500 126.800 ;
        RECT 18.200 126.200 18.500 126.800 ;
        RECT 23.800 126.200 24.100 127.800 ;
        RECT 27.000 127.200 27.300 127.800 ;
        RECT 27.800 127.200 28.100 127.800 ;
        RECT 31.800 127.200 32.100 127.800 ;
        RECT 27.000 126.800 27.400 127.200 ;
        RECT 27.800 126.800 28.200 127.200 ;
        RECT 31.800 126.800 32.200 127.200 ;
        RECT 34.200 126.800 34.600 127.200 ;
        RECT 11.000 126.100 11.400 126.200 ;
        RECT 11.800 126.100 12.200 126.200 ;
        RECT 11.000 125.800 12.200 126.100 ;
        RECT 14.200 125.800 14.600 126.200 ;
        RECT 15.800 125.800 16.200 126.200 ;
        RECT 18.200 125.800 18.600 126.200 ;
        RECT 19.800 126.100 20.200 126.200 ;
        RECT 20.600 126.100 21.000 126.200 ;
        RECT 19.800 125.800 21.000 126.100 ;
        RECT 23.800 125.800 24.200 126.200 ;
        RECT 26.200 125.800 26.600 126.200 ;
        RECT 15.800 125.200 16.100 125.800 ;
        RECT 26.200 125.200 26.500 125.800 ;
        RECT 8.600 124.800 9.000 125.200 ;
        RECT 9.400 125.100 9.800 125.200 ;
        RECT 10.200 125.100 10.600 125.200 ;
        RECT 9.400 124.800 10.600 125.100 ;
        RECT 12.600 125.100 13.000 125.200 ;
        RECT 13.400 125.100 13.800 125.200 ;
        RECT 12.600 124.800 13.800 125.100 ;
        RECT 15.800 124.800 16.200 125.200 ;
        RECT 17.400 124.800 17.800 125.200 ;
        RECT 19.000 125.100 19.400 125.200 ;
        RECT 19.000 124.800 20.100 125.100 ;
        RECT 17.400 124.200 17.700 124.800 ;
        RECT 9.400 123.800 9.800 124.200 ;
        RECT 11.800 124.100 12.200 124.200 ;
        RECT 12.600 124.100 13.000 124.200 ;
        RECT 11.800 123.800 13.000 124.100 ;
        RECT 17.400 123.800 17.800 124.200 ;
        RECT 7.000 121.800 7.400 122.200 ;
        RECT 3.000 120.800 3.400 121.200 ;
        RECT 6.200 120.800 6.600 121.200 ;
        RECT 2.200 118.800 2.600 119.200 ;
        RECT 7.000 118.200 7.300 121.800 ;
        RECT 9.400 119.200 9.700 123.800 ;
        RECT 17.400 122.800 17.800 123.200 ;
        RECT 17.400 119.200 17.700 122.800 ;
        RECT 18.200 122.100 18.600 122.200 ;
        RECT 19.000 122.100 19.400 122.200 ;
        RECT 18.200 121.800 19.400 122.100 ;
        RECT 19.800 119.200 20.100 124.800 ;
        RECT 23.800 124.800 24.200 125.200 ;
        RECT 26.200 124.800 26.600 125.200 ;
        RECT 22.200 124.100 22.600 124.200 ;
        RECT 23.000 124.100 23.400 124.200 ;
        RECT 22.200 123.800 23.400 124.100 ;
        RECT 20.600 121.800 21.000 122.200 ;
        RECT 9.400 118.800 9.800 119.200 ;
        RECT 17.400 118.800 17.800 119.200 ;
        RECT 19.800 118.800 20.200 119.200 ;
        RECT 7.000 117.800 7.400 118.200 ;
        RECT 1.400 117.100 1.800 117.200 ;
        RECT 2.200 117.100 2.600 117.200 ;
        RECT 1.400 116.800 2.600 117.100 ;
        RECT 3.800 117.100 4.200 117.200 ;
        RECT 4.600 117.100 5.000 117.200 ;
        RECT 3.800 116.800 5.000 117.100 ;
        RECT 11.800 117.100 12.200 117.200 ;
        RECT 12.600 117.100 13.000 117.200 ;
        RECT 11.800 116.800 13.000 117.100 ;
        RECT 15.000 117.100 15.400 117.200 ;
        RECT 15.800 117.100 16.200 117.200 ;
        RECT 15.000 116.800 16.200 117.100 ;
        RECT 16.600 116.800 17.000 117.200 ;
        RECT 3.000 115.800 3.400 116.200 ;
        RECT 6.200 115.800 6.600 116.200 ;
        RECT 10.200 115.800 10.600 116.200 ;
        RECT 11.000 115.800 11.400 116.200 ;
        RECT 11.800 116.100 12.200 116.200 ;
        RECT 12.600 116.100 13.000 116.200 ;
        RECT 11.800 115.800 13.000 116.100 ;
        RECT 14.200 115.800 14.600 116.200 ;
        RECT 2.200 114.800 2.600 115.200 ;
        RECT 2.200 114.200 2.500 114.800 ;
        RECT 3.000 114.200 3.300 115.800 ;
        RECT 3.800 115.100 4.200 115.200 ;
        RECT 4.600 115.100 5.000 115.200 ;
        RECT 3.800 114.800 5.000 115.100 ;
        RECT 5.400 114.800 5.800 115.200 ;
        RECT 2.200 113.800 2.600 114.200 ;
        RECT 3.000 113.800 3.400 114.200 ;
        RECT 5.400 113.200 5.700 114.800 ;
        RECT 5.400 112.800 5.800 113.200 ;
        RECT 3.800 107.800 4.200 108.200 ;
        RECT 5.400 107.800 5.800 108.200 ;
        RECT 3.800 107.200 4.100 107.800 ;
        RECT 5.400 107.200 5.700 107.800 ;
        RECT 3.800 106.800 4.200 107.200 ;
        RECT 5.400 106.800 5.800 107.200 ;
        RECT 6.200 106.200 6.500 115.800 ;
        RECT 7.000 114.800 7.400 115.200 ;
        RECT 7.000 114.200 7.300 114.800 ;
        RECT 7.000 113.800 7.400 114.200 ;
        RECT 8.600 112.800 9.000 113.200 ;
        RECT 7.800 111.800 8.200 112.200 ;
        RECT 7.800 106.200 8.100 111.800 ;
        RECT 8.600 109.200 8.900 112.800 ;
        RECT 8.600 108.800 9.000 109.200 ;
        RECT 8.600 106.800 9.000 107.200 ;
        RECT 8.600 106.200 8.900 106.800 ;
        RECT 3.000 106.100 3.400 106.200 ;
        RECT 3.800 106.100 4.200 106.200 ;
        RECT 3.000 105.800 4.200 106.100 ;
        RECT 6.200 105.800 6.600 106.200 ;
        RECT 7.800 105.800 8.200 106.200 ;
        RECT 8.600 105.800 9.000 106.200 ;
        RECT 6.200 105.200 6.500 105.800 ;
        RECT 0.600 105.100 1.000 105.200 ;
        RECT 1.400 105.100 1.800 105.200 ;
        RECT 0.600 104.800 1.800 105.100 ;
        RECT 2.200 104.800 2.600 105.200 ;
        RECT 6.200 104.800 6.600 105.200 ;
        RECT 8.600 105.100 9.000 105.200 ;
        RECT 9.400 105.100 9.800 105.200 ;
        RECT 8.600 104.800 9.800 105.100 ;
        RECT 2.200 104.200 2.500 104.800 ;
        RECT 2.200 103.800 2.600 104.200 ;
        RECT 2.200 101.800 2.600 102.200 ;
        RECT 8.600 101.800 9.000 102.200 ;
        RECT 2.200 99.200 2.500 101.800 ;
        RECT 2.200 98.800 2.600 99.200 ;
        RECT 7.000 99.100 7.400 99.200 ;
        RECT 7.800 99.100 8.200 99.200 ;
        RECT 7.000 98.800 8.200 99.100 ;
        RECT 8.600 97.200 8.900 101.800 ;
        RECT 10.200 99.200 10.500 115.800 ;
        RECT 11.000 115.200 11.300 115.800 ;
        RECT 11.000 114.800 11.400 115.200 ;
        RECT 11.000 113.200 11.300 114.800 ;
        RECT 14.200 114.200 14.500 115.800 ;
        RECT 16.600 115.200 16.900 116.800 ;
        RECT 18.200 116.100 18.600 116.200 ;
        RECT 18.200 115.800 19.300 116.100 ;
        RECT 15.000 114.800 15.400 115.200 ;
        RECT 16.600 114.800 17.000 115.200 ;
        RECT 14.200 113.800 14.600 114.200 ;
        RECT 11.000 112.800 11.400 113.200 ;
        RECT 12.600 111.800 13.000 112.200 ;
        RECT 11.000 108.800 11.400 109.200 ;
        RECT 11.000 106.200 11.300 108.800 ;
        RECT 12.600 108.200 12.900 111.800 ;
        RECT 12.600 107.800 13.000 108.200 ;
        RECT 11.000 105.800 11.400 106.200 ;
        RECT 11.800 104.100 12.200 104.200 ;
        RECT 12.600 104.100 12.900 107.800 ;
        RECT 13.400 107.100 13.800 107.200 ;
        RECT 14.200 107.100 14.600 107.200 ;
        RECT 13.400 106.800 14.600 107.100 ;
        RECT 15.000 105.200 15.300 114.800 ;
        RECT 16.600 114.200 16.900 114.800 ;
        RECT 16.600 113.800 17.000 114.200 ;
        RECT 17.400 113.100 17.800 113.200 ;
        RECT 18.200 113.100 18.600 113.200 ;
        RECT 17.400 112.800 18.600 113.100 ;
        RECT 19.000 112.200 19.300 115.800 ;
        RECT 19.000 111.800 19.400 112.200 ;
        RECT 16.600 108.800 17.000 109.200 ;
        RECT 16.600 108.200 16.900 108.800 ;
        RECT 19.800 108.200 20.100 118.800 ;
        RECT 20.600 116.200 20.900 121.800 ;
        RECT 20.600 115.800 21.000 116.200 ;
        RECT 22.200 115.800 22.600 116.200 ;
        RECT 20.600 113.800 21.000 114.200 ;
        RECT 21.400 113.800 21.800 114.200 ;
        RECT 20.600 111.200 20.900 113.800 ;
        RECT 21.400 113.200 21.700 113.800 ;
        RECT 21.400 112.800 21.800 113.200 ;
        RECT 20.600 110.800 21.000 111.200 ;
        RECT 16.600 107.800 17.000 108.200 ;
        RECT 19.800 107.800 20.200 108.200 ;
        RECT 15.800 107.100 16.200 107.200 ;
        RECT 16.600 107.100 17.000 107.200 ;
        RECT 15.800 106.800 17.000 107.100 ;
        RECT 17.400 105.800 17.800 106.200 ;
        RECT 20.600 106.100 21.000 106.200 ;
        RECT 21.400 106.100 21.800 106.200 ;
        RECT 20.600 105.800 21.800 106.100 ;
        RECT 15.000 104.800 15.400 105.200 ;
        RECT 11.800 103.800 12.900 104.100 ;
        RECT 12.600 101.800 13.000 102.200 ;
        RECT 14.200 101.800 14.600 102.200 ;
        RECT 10.200 98.800 10.600 99.200 ;
        RECT 1.400 97.100 1.800 97.200 ;
        RECT 2.200 97.100 2.600 97.200 ;
        RECT 1.400 96.800 2.600 97.100 ;
        RECT 5.400 97.100 5.800 97.200 ;
        RECT 6.200 97.100 6.600 97.200 ;
        RECT 5.400 96.800 6.600 97.100 ;
        RECT 8.600 96.800 9.000 97.200 ;
        RECT 3.000 95.800 3.400 96.200 ;
        RECT 7.800 95.800 8.200 96.200 ;
        RECT 8.600 96.100 9.000 96.200 ;
        RECT 9.400 96.100 9.800 96.200 ;
        RECT 8.600 95.800 9.800 96.100 ;
        RECT 1.400 94.800 1.800 95.200 ;
        RECT 0.600 93.800 1.000 94.200 ;
        RECT 0.600 86.200 0.900 93.800 ;
        RECT 1.400 89.200 1.700 94.800 ;
        RECT 3.000 94.200 3.300 95.800 ;
        RECT 4.600 94.800 5.000 95.200 ;
        RECT 6.200 95.100 6.600 95.200 ;
        RECT 7.000 95.100 7.400 95.200 ;
        RECT 6.200 94.800 7.400 95.100 ;
        RECT 3.000 94.100 3.400 94.200 ;
        RECT 3.800 94.100 4.200 94.200 ;
        RECT 3.000 93.800 4.200 94.100 ;
        RECT 2.200 92.800 2.600 93.200 ;
        RECT 1.400 88.800 1.800 89.200 ;
        RECT 1.400 87.200 1.700 88.800 ;
        RECT 1.400 86.800 1.800 87.200 ;
        RECT 0.600 85.800 1.000 86.200 ;
        RECT 0.600 85.200 0.900 85.800 ;
        RECT 0.600 84.800 1.000 85.200 ;
        RECT 2.200 79.200 2.500 92.800 ;
        RECT 4.600 92.200 4.900 94.800 ;
        RECT 3.800 91.800 4.200 92.200 ;
        RECT 4.600 91.800 5.000 92.200 ;
        RECT 3.800 89.200 4.100 91.800 ;
        RECT 3.800 88.800 4.200 89.200 ;
        RECT 3.000 87.800 3.400 88.200 ;
        RECT 4.600 88.100 4.900 91.800 ;
        RECT 7.800 89.200 8.100 95.800 ;
        RECT 11.000 94.800 11.400 95.200 ;
        RECT 12.600 95.100 12.900 101.800 ;
        RECT 14.200 95.200 14.500 101.800 ;
        RECT 17.400 101.100 17.700 105.800 ;
        RECT 22.200 105.200 22.500 115.800 ;
        RECT 23.800 115.200 24.100 124.800 ;
        RECT 24.600 124.100 25.000 124.200 ;
        RECT 25.400 124.100 25.800 124.200 ;
        RECT 24.600 123.800 25.800 124.100 ;
        RECT 27.000 123.200 27.300 126.800 ;
        RECT 29.400 125.800 29.800 126.200 ;
        RECT 30.200 126.100 30.600 126.200 ;
        RECT 31.000 126.100 31.400 126.200 ;
        RECT 30.200 125.800 31.400 126.100 ;
        RECT 29.400 123.200 29.700 125.800 ;
        RECT 27.000 122.800 27.400 123.200 ;
        RECT 29.400 122.800 29.800 123.200 ;
        RECT 31.800 119.200 32.100 126.800 ;
        RECT 31.800 118.800 32.200 119.200 ;
        RECT 27.000 117.800 27.400 118.200 ;
        RECT 27.000 117.200 27.300 117.800 ;
        RECT 25.400 116.800 25.800 117.200 ;
        RECT 27.000 116.800 27.400 117.200 ;
        RECT 25.400 116.200 25.700 116.800 ;
        RECT 25.400 115.800 25.800 116.200 ;
        RECT 28.600 115.800 29.000 116.200 ;
        RECT 30.200 115.800 30.600 116.200 ;
        RECT 23.000 114.800 23.400 115.200 ;
        RECT 23.800 114.800 24.200 115.200 ;
        RECT 26.200 115.100 26.600 115.200 ;
        RECT 25.400 114.800 26.600 115.100 ;
        RECT 23.000 114.200 23.300 114.800 ;
        RECT 23.000 113.800 23.400 114.200 ;
        RECT 23.800 113.800 24.200 114.200 ;
        RECT 23.000 110.200 23.300 113.800 ;
        RECT 23.800 113.200 24.100 113.800 ;
        RECT 25.400 113.200 25.700 114.800 ;
        RECT 28.600 114.200 28.900 115.800 ;
        RECT 29.400 114.800 29.800 115.200 ;
        RECT 26.200 114.100 26.600 114.200 ;
        RECT 26.200 113.800 27.300 114.100 ;
        RECT 23.800 112.800 24.200 113.200 ;
        RECT 25.400 112.800 25.800 113.200 ;
        RECT 23.000 109.800 23.400 110.200 ;
        RECT 25.400 109.200 25.700 112.800 ;
        RECT 27.000 111.200 27.300 113.800 ;
        RECT 28.600 113.800 29.000 114.200 ;
        RECT 27.000 110.800 27.400 111.200 ;
        RECT 27.000 109.200 27.300 110.800 ;
        RECT 25.400 108.800 25.800 109.200 ;
        RECT 27.000 108.800 27.400 109.200 ;
        RECT 28.600 108.200 28.900 113.800 ;
        RECT 29.400 113.200 29.700 114.800 ;
        RECT 30.200 114.200 30.500 115.800 ;
        RECT 31.800 114.200 32.100 118.800 ;
        RECT 34.200 118.200 34.500 126.800 ;
        RECT 40.600 126.200 40.900 127.800 ;
        RECT 41.400 127.100 41.800 127.200 ;
        RECT 42.200 127.100 42.600 127.200 ;
        RECT 41.400 126.800 42.600 127.100 ;
        RECT 45.400 127.100 45.800 127.200 ;
        RECT 46.200 127.100 46.600 127.200 ;
        RECT 45.400 126.800 46.600 127.100 ;
        RECT 35.000 126.100 35.400 126.200 ;
        RECT 35.800 126.100 36.200 126.200 ;
        RECT 35.000 125.800 36.200 126.100 ;
        RECT 39.800 125.800 40.200 126.200 ;
        RECT 40.600 125.800 41.000 126.200 ;
        RECT 42.200 126.100 42.600 126.200 ;
        RECT 43.000 126.100 43.400 126.200 ;
        RECT 42.200 125.800 43.400 126.100 ;
        RECT 45.400 125.800 45.800 126.200 ;
        RECT 36.600 124.900 37.000 125.300 ;
        RECT 38.200 125.100 38.600 125.200 ;
        RECT 39.000 125.100 39.400 125.200 ;
        RECT 36.600 124.200 36.900 124.900 ;
        RECT 38.200 124.800 39.400 125.100 ;
        RECT 36.600 123.800 37.000 124.200 ;
        RECT 38.200 123.800 38.600 124.200 ;
        RECT 35.800 122.800 36.200 123.200 ;
        RECT 34.200 117.800 34.600 118.200 ;
        RECT 33.400 116.800 33.800 117.200 ;
        RECT 33.400 116.200 33.700 116.800 ;
        RECT 35.800 116.200 36.100 122.800 ;
        RECT 38.200 121.200 38.500 123.800 ;
        RECT 38.200 120.800 38.600 121.200 ;
        RECT 38.200 119.200 38.500 120.800 ;
        RECT 38.200 118.800 38.600 119.200 ;
        RECT 39.000 117.800 39.400 118.200 ;
        RECT 36.600 117.100 37.000 117.200 ;
        RECT 37.400 117.100 37.800 117.200 ;
        RECT 36.600 116.800 37.800 117.100 ;
        RECT 39.000 116.200 39.300 117.800 ;
        RECT 33.400 115.800 33.800 116.200 ;
        RECT 35.000 115.800 35.400 116.200 ;
        RECT 35.800 115.800 36.200 116.200 ;
        RECT 39.000 115.800 39.400 116.200 ;
        RECT 33.400 114.800 33.800 115.200 ;
        RECT 34.200 114.800 34.600 115.200 ;
        RECT 33.400 114.200 33.700 114.800 ;
        RECT 30.200 113.800 30.600 114.200 ;
        RECT 31.800 113.800 32.200 114.200 ;
        RECT 33.400 113.800 33.800 114.200 ;
        RECT 29.400 112.800 29.800 113.200 ;
        RECT 30.200 112.200 30.500 113.800 ;
        RECT 34.200 113.200 34.500 114.800 ;
        RECT 31.800 112.800 32.200 113.200 ;
        RECT 34.200 112.800 34.600 113.200 ;
        RECT 30.200 111.800 30.600 112.200 ;
        RECT 30.200 109.200 30.500 111.800 ;
        RECT 31.800 111.200 32.100 112.800 ;
        RECT 34.200 112.200 34.500 112.800 ;
        RECT 34.200 111.800 34.600 112.200 ;
        RECT 35.000 111.200 35.300 115.800 ;
        RECT 35.800 115.100 36.200 115.200 ;
        RECT 36.600 115.100 37.000 115.200 ;
        RECT 35.800 114.800 37.000 115.100 ;
        RECT 39.800 115.100 40.100 125.800 ;
        RECT 41.400 124.800 41.800 125.200 ;
        RECT 44.600 124.800 45.000 125.200 ;
        RECT 41.400 124.200 41.700 124.800 ;
        RECT 40.600 123.800 41.000 124.200 ;
        RECT 41.400 123.800 41.800 124.200 ;
        RECT 40.600 119.200 40.900 123.800 ;
        RECT 44.600 123.200 44.900 124.800 ;
        RECT 44.600 122.800 45.000 123.200 ;
        RECT 45.400 122.100 45.700 125.800 ;
        RECT 47.800 124.200 48.100 127.800 ;
        RECT 51.000 126.800 51.400 127.200 ;
        RECT 59.800 126.800 60.200 127.200 ;
        RECT 51.000 126.200 51.300 126.800 ;
        RECT 59.800 126.200 60.100 126.800 ;
        RECT 61.400 126.200 61.700 127.800 ;
        RECT 62.200 126.200 62.500 127.800 ;
        RECT 63.000 127.100 63.400 127.200 ;
        RECT 63.800 127.100 64.200 127.200 ;
        RECT 63.000 126.800 64.200 127.100 ;
        RECT 64.600 127.100 65.000 127.200 ;
        RECT 65.400 127.100 65.800 127.200 ;
        RECT 64.600 126.800 65.800 127.100 ;
        RECT 66.200 127.100 66.600 127.200 ;
        RECT 67.000 127.100 67.400 127.200 ;
        RECT 66.200 126.800 67.400 127.100 ;
        RECT 68.600 126.800 69.000 127.200 ;
        RECT 68.600 126.200 68.900 126.800 ;
        RECT 71.800 126.200 72.100 127.800 ;
        RECT 74.200 126.800 74.600 127.200 ;
        RECT 77.400 127.100 77.800 127.200 ;
        RECT 78.200 127.100 78.600 127.200 ;
        RECT 77.400 126.800 78.600 127.100 ;
        RECT 84.600 126.800 85.000 127.200 ;
        RECT 74.200 126.200 74.500 126.800 ;
        RECT 84.600 126.200 84.900 126.800 ;
        RECT 50.200 125.800 50.600 126.200 ;
        RECT 51.000 125.800 51.400 126.200 ;
        RECT 55.000 125.800 55.400 126.200 ;
        RECT 59.800 125.800 60.200 126.200 ;
        RECT 61.400 125.800 61.800 126.200 ;
        RECT 62.200 125.800 62.600 126.200 ;
        RECT 65.400 125.800 65.800 126.200 ;
        RECT 68.600 125.800 69.000 126.200 ;
        RECT 71.800 125.800 72.200 126.200 ;
        RECT 74.200 125.800 74.600 126.200 ;
        RECT 75.800 125.800 76.200 126.200 ;
        RECT 80.600 126.100 81.000 126.200 ;
        RECT 81.400 126.100 81.800 126.200 ;
        RECT 80.600 125.800 81.800 126.100 ;
        RECT 84.600 125.800 85.000 126.200 ;
        RECT 50.200 125.200 50.500 125.800 ;
        RECT 55.000 125.200 55.300 125.800 ;
        RECT 50.200 124.800 50.600 125.200 ;
        RECT 55.000 124.800 55.400 125.200 ;
        RECT 55.800 124.800 56.200 125.200 ;
        RECT 47.800 123.800 48.200 124.200 ;
        RECT 51.000 124.100 51.400 124.200 ;
        RECT 51.800 124.100 52.200 124.200 ;
        RECT 51.000 123.800 52.200 124.100 ;
        RECT 52.600 124.100 53.000 124.200 ;
        RECT 54.200 124.100 54.600 124.200 ;
        RECT 52.600 123.800 54.600 124.100 ;
        RECT 44.600 121.800 45.700 122.100 ;
        RECT 55.000 121.800 55.400 122.200 ;
        RECT 44.600 119.200 44.900 121.800 ;
        RECT 55.000 121.200 55.300 121.800 ;
        RECT 55.000 120.800 55.400 121.200 ;
        RECT 55.000 119.800 55.400 120.200 ;
        RECT 55.000 119.200 55.300 119.800 ;
        RECT 55.800 119.200 56.100 124.800 ;
        RECT 59.800 123.200 60.100 125.800 ;
        RECT 59.800 122.800 60.200 123.200 ;
        RECT 59.800 120.200 60.100 122.800 ;
        RECT 59.800 119.800 60.200 120.200 ;
        RECT 40.600 118.800 41.000 119.200 ;
        RECT 44.600 118.800 45.000 119.200 ;
        RECT 55.000 118.800 55.400 119.200 ;
        RECT 55.800 118.800 56.200 119.200 ;
        RECT 59.000 118.800 59.400 119.200 ;
        RECT 59.000 118.200 59.300 118.800 ;
        RECT 42.200 117.800 42.600 118.200 ;
        RECT 59.000 117.800 59.400 118.200 ;
        RECT 42.200 116.200 42.500 117.800 ;
        RECT 43.000 117.100 43.400 117.200 ;
        RECT 43.800 117.100 44.200 117.200 ;
        RECT 43.000 116.800 44.200 117.100 ;
        RECT 42.200 115.800 42.600 116.200 ;
        RECT 53.400 115.800 53.800 116.200 ;
        RECT 40.600 115.100 41.000 115.200 ;
        RECT 39.800 114.800 41.000 115.100 ;
        RECT 42.200 115.100 42.600 115.200 ;
        RECT 43.000 115.100 43.400 115.200 ;
        RECT 42.200 114.800 43.400 115.100 ;
        RECT 39.800 113.200 40.100 114.800 ;
        RECT 40.600 114.100 41.000 114.200 ;
        RECT 41.400 114.100 41.800 114.200 ;
        RECT 40.600 113.800 41.800 114.100 ;
        RECT 47.000 113.800 47.400 114.200 ;
        RECT 51.800 113.800 52.200 114.200 ;
        RECT 36.600 112.800 37.000 113.200 ;
        RECT 39.800 112.800 40.200 113.200 ;
        RECT 45.400 112.800 45.800 113.200 ;
        RECT 31.800 110.800 32.200 111.200 ;
        RECT 35.000 110.800 35.400 111.200 ;
        RECT 36.600 109.200 36.900 112.800 ;
        RECT 45.400 112.200 45.700 112.800 ;
        RECT 43.000 111.800 43.400 112.200 ;
        RECT 45.400 111.800 45.800 112.200 ;
        RECT 46.200 111.800 46.600 112.200 ;
        RECT 43.000 109.200 43.300 111.800 ;
        RECT 30.200 108.800 30.600 109.200 ;
        RECT 36.600 108.800 37.000 109.200 ;
        RECT 39.800 109.100 40.200 109.200 ;
        RECT 40.600 109.100 41.000 109.200 ;
        RECT 39.800 108.800 41.000 109.100 ;
        RECT 43.000 108.800 43.400 109.200 ;
        RECT 24.600 107.800 25.000 108.200 ;
        RECT 25.400 107.800 25.800 108.200 ;
        RECT 26.200 107.800 26.600 108.200 ;
        RECT 28.600 107.800 29.000 108.200 ;
        RECT 35.000 108.100 35.400 108.200 ;
        RECT 35.800 108.100 36.200 108.200 ;
        RECT 35.000 107.800 36.200 108.100 ;
        RECT 39.000 107.800 39.400 108.200 ;
        RECT 24.600 107.200 24.900 107.800 ;
        RECT 24.600 106.800 25.000 107.200 ;
        RECT 25.400 106.200 25.700 107.800 ;
        RECT 24.600 105.800 25.000 106.200 ;
        RECT 25.400 105.800 25.800 106.200 ;
        RECT 18.200 105.100 18.600 105.200 ;
        RECT 19.000 105.100 19.400 105.200 ;
        RECT 18.200 104.800 19.400 105.100 ;
        RECT 22.200 104.800 22.600 105.200 ;
        RECT 19.800 104.100 20.200 104.200 ;
        RECT 20.600 104.100 21.000 104.200 ;
        RECT 19.800 103.800 21.000 104.100 ;
        RECT 21.400 103.800 21.800 104.200 ;
        RECT 23.000 104.100 23.400 104.200 ;
        RECT 23.800 104.100 24.200 104.200 ;
        RECT 23.000 103.800 24.200 104.100 ;
        RECT 21.400 103.200 21.700 103.800 ;
        RECT 24.600 103.200 24.900 105.800 ;
        RECT 26.200 104.200 26.500 107.800 ;
        RECT 39.000 107.200 39.300 107.800 ;
        RECT 46.200 107.200 46.500 111.800 ;
        RECT 47.000 107.200 47.300 113.800 ;
        RECT 51.000 112.800 51.400 113.200 ;
        RECT 50.200 111.800 50.600 112.200 ;
        RECT 27.800 106.800 28.200 107.200 ;
        RECT 34.200 106.800 34.600 107.200 ;
        RECT 37.400 106.800 37.800 107.200 ;
        RECT 39.000 106.800 39.400 107.200 ;
        RECT 40.600 106.800 41.000 107.200 ;
        RECT 43.800 106.800 44.200 107.200 ;
        RECT 46.200 106.800 46.600 107.200 ;
        RECT 47.000 106.800 47.400 107.200 ;
        RECT 26.200 103.800 26.600 104.200 ;
        RECT 27.800 103.200 28.100 106.800 ;
        RECT 30.200 105.800 30.600 106.200 ;
        RECT 33.400 105.800 33.800 106.200 ;
        RECT 29.400 104.800 29.800 105.200 ;
        RECT 21.400 102.800 21.800 103.200 ;
        RECT 22.200 102.800 22.600 103.200 ;
        RECT 24.600 102.800 25.000 103.200 ;
        RECT 27.800 102.800 28.200 103.200 ;
        RECT 16.600 100.800 17.700 101.100 ;
        RECT 18.200 101.800 18.600 102.200 ;
        RECT 16.600 99.200 16.900 100.800 ;
        RECT 16.600 98.800 17.000 99.200 ;
        RECT 15.800 96.800 16.200 97.200 ;
        RECT 16.600 96.800 17.000 97.200 ;
        RECT 15.800 96.200 16.100 96.800 ;
        RECT 15.800 95.800 16.200 96.200 ;
        RECT 16.600 95.200 16.900 96.800 ;
        RECT 17.400 96.100 17.800 96.200 ;
        RECT 18.200 96.100 18.500 101.800 ;
        RECT 22.200 99.200 22.500 102.800 ;
        RECT 29.400 99.200 29.700 104.800 ;
        RECT 30.200 103.200 30.500 105.800 ;
        RECT 31.800 105.100 32.200 105.200 ;
        RECT 32.600 105.100 33.000 105.200 ;
        RECT 31.800 104.800 33.000 105.100 ;
        RECT 31.000 104.100 31.400 104.200 ;
        RECT 31.800 104.100 32.200 104.200 ;
        RECT 31.000 103.800 32.200 104.100 ;
        RECT 32.600 103.800 33.000 104.200 ;
        RECT 30.200 102.800 30.600 103.200 ;
        RECT 32.600 99.200 32.900 103.800 ;
        RECT 33.400 103.200 33.700 105.800 ;
        RECT 34.200 104.200 34.500 106.800 ;
        RECT 37.400 106.200 37.700 106.800 ;
        RECT 40.600 106.200 40.900 106.800 ;
        RECT 35.000 105.800 35.400 106.200 ;
        RECT 37.400 105.800 37.800 106.200 ;
        RECT 38.200 105.800 38.600 106.200 ;
        RECT 40.600 105.800 41.000 106.200 ;
        RECT 42.200 106.100 42.600 106.200 ;
        RECT 43.000 106.100 43.400 106.200 ;
        RECT 42.200 105.800 43.400 106.100 ;
        RECT 35.000 105.200 35.300 105.800 ;
        RECT 38.200 105.200 38.500 105.800 ;
        RECT 35.000 104.800 35.400 105.200 ;
        RECT 38.200 104.800 38.600 105.200 ;
        RECT 40.600 104.200 40.900 105.800 ;
        RECT 42.200 105.100 42.600 105.200 ;
        RECT 43.000 105.100 43.400 105.200 ;
        RECT 42.200 104.800 43.400 105.100 ;
        RECT 43.800 104.200 44.100 106.800 ;
        RECT 45.400 106.100 45.800 106.200 ;
        RECT 46.200 106.100 46.600 106.200 ;
        RECT 45.400 105.800 46.600 106.100 ;
        RECT 47.800 106.100 48.200 106.200 ;
        RECT 48.600 106.100 49.000 106.200 ;
        RECT 47.800 105.800 49.000 106.100 ;
        RECT 50.200 105.200 50.500 111.800 ;
        RECT 51.000 108.200 51.300 112.800 ;
        RECT 51.800 109.200 52.100 113.800 ;
        RECT 51.800 108.800 52.200 109.200 ;
        RECT 51.000 107.800 51.400 108.200 ;
        RECT 51.000 106.800 51.400 107.200 ;
        RECT 51.000 106.200 51.300 106.800 ;
        RECT 53.400 106.200 53.700 115.800 ;
        RECT 61.400 114.800 61.800 115.200 ;
        RECT 61.400 114.200 61.700 114.800 ;
        RECT 54.200 113.800 54.600 114.200 ;
        RECT 57.400 114.100 57.800 114.200 ;
        RECT 58.200 114.100 58.600 114.200 ;
        RECT 57.400 113.800 58.600 114.100 ;
        RECT 59.800 114.100 60.200 114.200 ;
        RECT 60.600 114.100 61.000 114.200 ;
        RECT 59.800 113.800 61.000 114.100 ;
        RECT 61.400 113.800 61.800 114.200 ;
        RECT 54.200 113.200 54.500 113.800 ;
        RECT 54.200 112.800 54.600 113.200 ;
        RECT 55.800 113.100 56.200 113.200 ;
        RECT 56.600 113.100 57.000 113.200 ;
        RECT 55.800 112.800 57.000 113.100 ;
        RECT 59.800 112.800 60.200 113.200 ;
        RECT 62.200 113.100 62.500 125.800 ;
        RECT 65.400 125.200 65.700 125.800 ;
        RECT 65.400 124.800 65.800 125.200 ;
        RECT 67.800 124.800 68.200 125.200 ;
        RECT 71.000 125.100 71.400 125.200 ;
        RECT 69.400 124.800 71.400 125.100 ;
        RECT 73.400 125.100 73.800 125.200 ;
        RECT 74.200 125.100 74.600 125.200 ;
        RECT 73.400 124.800 74.600 125.100 ;
        RECT 64.600 119.800 65.000 120.200 ;
        RECT 64.600 119.200 64.900 119.800 ;
        RECT 67.800 119.200 68.100 124.800 ;
        RECT 69.400 124.200 69.700 124.800 ;
        RECT 69.400 123.800 69.800 124.200 ;
        RECT 70.200 123.800 70.600 124.200 ;
        RECT 72.600 124.100 73.000 124.200 ;
        RECT 73.400 124.100 73.800 124.200 ;
        RECT 72.600 123.800 73.800 124.100 ;
        RECT 70.200 123.200 70.500 123.800 ;
        RECT 70.200 122.800 70.600 123.200 ;
        RECT 74.200 121.800 74.600 122.200 ;
        RECT 74.200 119.200 74.500 121.800 ;
        RECT 75.800 119.200 76.100 125.800 ;
        RECT 81.400 125.100 81.800 125.200 ;
        RECT 82.200 125.100 82.600 125.200 ;
        RECT 81.400 124.800 82.600 125.100 ;
        RECT 80.600 123.800 81.000 124.200 ;
        RECT 79.000 119.800 79.400 120.200 ;
        RECT 64.600 118.800 65.000 119.200 ;
        RECT 67.800 118.800 68.200 119.200 ;
        RECT 74.200 118.800 74.600 119.200 ;
        RECT 75.800 118.800 76.200 119.200 ;
        RECT 71.800 117.800 72.200 118.200 ;
        RECT 71.800 117.200 72.100 117.800 ;
        RECT 69.400 116.800 69.800 117.200 ;
        RECT 71.800 116.800 72.200 117.200 ;
        RECT 74.200 117.100 74.600 117.200 ;
        RECT 75.000 117.100 75.400 117.200 ;
        RECT 74.200 116.800 75.400 117.100 ;
        RECT 61.400 112.800 62.500 113.100 ;
        RECT 63.000 115.800 63.400 116.200 ;
        RECT 67.000 116.100 67.400 116.200 ;
        RECT 67.800 116.100 68.200 116.200 ;
        RECT 67.000 115.800 68.200 116.100 ;
        RECT 63.000 114.200 63.300 115.800 ;
        RECT 66.200 114.800 66.600 115.200 ;
        RECT 67.000 114.800 67.400 115.200 ;
        RECT 67.800 115.100 68.200 115.200 ;
        RECT 68.600 115.100 69.000 115.200 ;
        RECT 67.800 114.800 69.000 115.100 ;
        RECT 66.200 114.200 66.500 114.800 ;
        RECT 63.000 113.800 63.400 114.200 ;
        RECT 63.800 114.100 64.200 114.200 ;
        RECT 64.600 114.100 65.000 114.200 ;
        RECT 63.800 113.800 65.000 114.100 ;
        RECT 66.200 113.800 66.600 114.200 ;
        RECT 63.000 113.200 63.300 113.800 ;
        RECT 66.200 113.200 66.500 113.800 ;
        RECT 63.000 112.800 63.400 113.200 ;
        RECT 63.800 113.100 64.200 113.200 ;
        RECT 64.600 113.100 65.000 113.200 ;
        RECT 63.800 112.800 65.000 113.100 ;
        RECT 66.200 112.800 66.600 113.200 ;
        RECT 59.800 112.200 60.100 112.800 ;
        RECT 59.800 111.800 60.200 112.200 ;
        RECT 56.600 110.800 57.000 111.200 ;
        RECT 55.000 107.800 55.400 108.200 ;
        RECT 55.000 106.200 55.300 107.800 ;
        RECT 55.800 106.800 56.200 107.200 ;
        RECT 51.000 105.800 51.400 106.200 ;
        RECT 53.400 105.800 53.800 106.200 ;
        RECT 55.000 105.800 55.400 106.200 ;
        RECT 45.400 104.800 45.800 105.200 ;
        RECT 50.200 104.800 50.600 105.200 ;
        RECT 34.200 103.800 34.600 104.200 ;
        RECT 40.600 103.800 41.000 104.200 ;
        RECT 43.800 103.800 44.200 104.200 ;
        RECT 33.400 102.800 33.800 103.200 ;
        RECT 45.400 99.200 45.700 104.800 ;
        RECT 47.000 104.100 47.400 104.200 ;
        RECT 47.800 104.100 48.200 104.200 ;
        RECT 47.000 103.800 48.200 104.100 ;
        RECT 46.200 102.800 46.600 103.200 ;
        RECT 46.200 99.200 46.500 102.800 ;
        RECT 51.000 101.200 51.300 105.800 ;
        RECT 53.400 104.800 53.800 105.200 ;
        RECT 55.000 104.800 55.400 105.200 ;
        RECT 51.800 103.800 52.200 104.200 ;
        RECT 51.800 103.200 52.100 103.800 ;
        RECT 53.400 103.200 53.700 104.800 ;
        RECT 55.000 104.200 55.300 104.800 ;
        RECT 55.000 103.800 55.400 104.200 ;
        RECT 51.800 102.800 52.200 103.200 ;
        RECT 53.400 102.800 53.800 103.200 ;
        RECT 55.800 102.200 56.100 106.800 ;
        RECT 55.800 101.800 56.200 102.200 ;
        RECT 51.000 100.800 51.400 101.200 ;
        RECT 56.600 99.200 56.900 110.800 ;
        RECT 61.400 109.200 61.700 112.800 ;
        RECT 60.600 108.800 61.000 109.200 ;
        RECT 61.400 108.800 61.800 109.200 ;
        RECT 62.200 108.800 62.600 109.200 ;
        RECT 66.200 108.800 66.600 109.200 ;
        RECT 60.600 107.200 60.900 108.800 ;
        RECT 62.200 108.200 62.500 108.800 ;
        RECT 66.200 108.200 66.500 108.800 ;
        RECT 62.200 107.800 62.600 108.200 ;
        RECT 64.600 107.800 65.000 108.200 ;
        RECT 66.200 107.800 66.600 108.200 ;
        RECT 64.600 107.200 64.900 107.800 ;
        RECT 58.200 107.100 58.600 107.200 ;
        RECT 59.000 107.100 59.400 107.200 ;
        RECT 58.200 106.800 59.400 107.100 ;
        RECT 60.600 106.800 61.000 107.200 ;
        RECT 63.000 106.800 63.400 107.200 ;
        RECT 64.600 106.800 65.000 107.200 ;
        RECT 63.000 106.200 63.300 106.800 ;
        RECT 57.400 106.100 57.800 106.200 ;
        RECT 58.200 106.100 58.600 106.200 ;
        RECT 57.400 105.800 58.600 106.100 ;
        RECT 59.000 105.800 59.400 106.200 ;
        RECT 59.800 105.800 60.200 106.200 ;
        RECT 63.000 105.800 63.400 106.200 ;
        RECT 63.800 105.800 64.200 106.200 ;
        RECT 59.000 104.200 59.300 105.800 ;
        RECT 59.800 105.200 60.100 105.800 ;
        RECT 59.800 104.800 60.200 105.200 ;
        RECT 59.000 103.800 59.400 104.200 ;
        RECT 62.200 103.800 62.600 104.200 ;
        RECT 59.000 100.800 59.400 101.200 ;
        RECT 59.000 99.200 59.300 100.800 ;
        RECT 62.200 99.200 62.500 103.800 ;
        RECT 22.200 98.800 22.600 99.200 ;
        RECT 29.400 98.800 29.800 99.200 ;
        RECT 32.600 98.800 33.000 99.200 ;
        RECT 45.400 98.800 45.800 99.200 ;
        RECT 46.200 98.800 46.600 99.200 ;
        RECT 51.000 99.100 51.400 99.200 ;
        RECT 51.800 99.100 52.200 99.200 ;
        RECT 51.000 98.800 52.200 99.100 ;
        RECT 56.600 98.800 57.000 99.200 ;
        RECT 59.000 98.800 59.400 99.200 ;
        RECT 62.200 98.800 62.600 99.200 ;
        RECT 26.200 97.800 26.600 98.200 ;
        RECT 28.600 97.800 29.000 98.200 ;
        RECT 31.800 97.800 32.200 98.200 ;
        RECT 38.200 97.800 38.600 98.200 ;
        RECT 40.600 97.800 41.000 98.200 ;
        RECT 47.000 97.800 47.400 98.200 ;
        RECT 51.800 97.800 52.200 98.200 ;
        RECT 54.200 97.800 54.600 98.200 ;
        RECT 17.400 95.800 18.500 96.100 ;
        RECT 18.200 95.200 18.500 95.800 ;
        RECT 19.000 96.800 19.400 97.200 ;
        RECT 12.600 94.800 13.700 95.100 ;
        RECT 14.200 94.800 14.600 95.200 ;
        RECT 16.600 94.800 17.000 95.200 ;
        RECT 18.200 94.800 18.600 95.200 ;
        RECT 8.600 93.800 9.000 94.200 ;
        RECT 8.600 93.200 8.900 93.800 ;
        RECT 8.600 92.800 9.000 93.200 ;
        RECT 10.200 91.800 10.600 92.200 ;
        RECT 7.000 89.100 7.400 89.200 ;
        RECT 7.800 89.100 8.200 89.200 ;
        RECT 7.000 88.800 8.200 89.100 ;
        RECT 10.200 88.200 10.500 91.800 ;
        RECT 3.800 87.800 4.900 88.100 ;
        RECT 7.800 87.800 8.200 88.200 ;
        RECT 10.200 87.800 10.600 88.200 ;
        RECT 3.000 86.200 3.300 87.800 ;
        RECT 3.000 85.800 3.400 86.200 ;
        RECT 3.800 85.200 4.100 87.800 ;
        RECT 6.200 87.100 6.600 87.200 ;
        RECT 7.000 87.100 7.400 87.200 ;
        RECT 6.200 86.800 7.400 87.100 ;
        RECT 4.600 86.100 5.000 86.200 ;
        RECT 5.400 86.100 5.800 86.200 ;
        RECT 4.600 85.800 5.800 86.100 ;
        RECT 3.800 84.800 4.200 85.200 ;
        RECT 3.000 81.800 3.400 82.200 ;
        RECT 2.200 78.800 2.600 79.200 ;
        RECT 1.400 76.800 1.800 77.200 ;
        RECT 1.400 67.200 1.700 76.800 ;
        RECT 3.000 76.200 3.300 81.800 ;
        RECT 3.800 79.200 4.100 84.800 ;
        RECT 7.800 84.200 8.100 87.800 ;
        RECT 8.600 86.800 9.000 87.200 ;
        RECT 8.600 86.200 8.900 86.800 ;
        RECT 8.600 85.800 9.000 86.200 ;
        RECT 9.400 86.100 9.800 86.200 ;
        RECT 10.200 86.100 10.600 86.200 ;
        RECT 9.400 85.800 10.600 86.100 ;
        RECT 9.400 84.800 9.800 85.200 ;
        RECT 7.800 83.800 8.200 84.200 ;
        RECT 8.600 83.800 9.000 84.200 ;
        RECT 7.800 79.200 8.100 83.800 ;
        RECT 3.800 78.800 4.200 79.200 ;
        RECT 5.400 78.800 5.800 79.200 ;
        RECT 7.800 78.800 8.200 79.200 ;
        RECT 3.000 75.800 3.400 76.200 ;
        RECT 3.800 75.800 4.200 76.200 ;
        RECT 2.200 74.800 2.600 75.200 ;
        RECT 1.400 66.800 1.800 67.200 ;
        RECT 0.600 65.800 1.000 66.200 ;
        RECT 0.600 65.200 0.900 65.800 ;
        RECT 0.600 64.800 1.000 65.200 ;
        RECT 0.600 52.800 1.000 53.200 ;
        RECT 0.600 52.200 0.900 52.800 ;
        RECT 0.600 51.800 1.000 52.200 ;
        RECT 1.400 45.100 1.700 66.800 ;
        RECT 2.200 65.200 2.500 74.800 ;
        RECT 3.000 68.200 3.300 75.800 ;
        RECT 3.800 75.200 4.100 75.800 ;
        RECT 5.400 75.200 5.700 78.800 ;
        RECT 7.800 76.800 8.200 77.200 ;
        RECT 6.200 76.100 6.600 76.200 ;
        RECT 7.000 76.100 7.400 76.200 ;
        RECT 6.200 75.800 7.400 76.100 ;
        RECT 3.800 74.800 4.200 75.200 ;
        RECT 5.400 74.800 5.800 75.200 ;
        RECT 6.200 74.800 6.600 75.200 ;
        RECT 6.200 74.200 6.500 74.800 ;
        RECT 7.800 74.200 8.100 76.800 ;
        RECT 8.600 75.200 8.900 83.800 ;
        RECT 9.400 82.200 9.700 84.800 ;
        RECT 9.400 81.800 9.800 82.200 ;
        RECT 9.400 76.100 9.800 76.200 ;
        RECT 10.200 76.100 10.600 76.200 ;
        RECT 9.400 75.800 10.600 76.100 ;
        RECT 8.600 74.800 9.000 75.200 ;
        RECT 9.400 75.100 9.800 75.200 ;
        RECT 10.200 75.100 10.600 75.200 ;
        RECT 9.400 74.800 10.600 75.100 ;
        RECT 4.600 73.800 5.000 74.200 ;
        RECT 6.200 73.800 6.600 74.200 ;
        RECT 7.800 73.800 8.200 74.200 ;
        RECT 4.600 70.100 4.900 73.800 ;
        RECT 8.600 73.200 8.900 74.800 ;
        RECT 8.600 72.800 9.000 73.200 ;
        RECT 9.400 73.100 9.800 73.200 ;
        RECT 10.200 73.100 10.600 73.200 ;
        RECT 9.400 72.800 10.600 73.100 ;
        RECT 4.600 69.800 5.700 70.100 ;
        RECT 4.600 68.800 5.000 69.200 ;
        RECT 4.600 68.200 4.900 68.800 ;
        RECT 5.400 68.200 5.700 69.800 ;
        RECT 11.000 69.200 11.300 94.800 ;
        RECT 13.400 94.200 13.700 94.800 ;
        RECT 19.000 94.200 19.300 96.800 ;
        RECT 20.600 95.800 21.000 96.200 ;
        RECT 23.000 96.100 23.400 96.200 ;
        RECT 23.800 96.100 24.200 96.200 ;
        RECT 23.000 95.800 24.200 96.100 ;
        RECT 11.800 93.800 12.200 94.200 ;
        RECT 12.600 93.800 13.000 94.200 ;
        RECT 13.400 93.800 13.800 94.200 ;
        RECT 19.000 93.800 19.400 94.200 ;
        RECT 11.800 93.200 12.100 93.800 ;
        RECT 12.600 93.200 12.900 93.800 ;
        RECT 20.600 93.200 20.900 95.800 ;
        RECT 22.200 94.800 22.600 95.200 ;
        RECT 22.200 94.200 22.500 94.800 ;
        RECT 26.200 94.200 26.500 97.800 ;
        RECT 28.600 97.200 28.900 97.800 ;
        RECT 31.800 97.200 32.100 97.800 ;
        RECT 38.200 97.200 38.500 97.800 ;
        RECT 40.600 97.200 40.900 97.800 ;
        RECT 47.000 97.200 47.300 97.800 ;
        RECT 51.800 97.200 52.100 97.800 ;
        RECT 54.200 97.200 54.500 97.800 ;
        RECT 28.600 96.800 29.000 97.200 ;
        RECT 31.800 96.800 32.200 97.200 ;
        RECT 34.200 96.800 34.600 97.200 ;
        RECT 38.200 96.800 38.600 97.200 ;
        RECT 39.000 97.100 39.400 97.200 ;
        RECT 39.800 97.100 40.200 97.200 ;
        RECT 39.000 96.800 40.200 97.100 ;
        RECT 40.600 96.800 41.000 97.200 ;
        RECT 43.000 97.100 43.400 97.200 ;
        RECT 43.800 97.100 44.200 97.200 ;
        RECT 43.000 96.800 44.200 97.100 ;
        RECT 46.200 96.800 46.600 97.200 ;
        RECT 47.000 96.800 47.400 97.200 ;
        RECT 51.000 96.800 51.400 97.200 ;
        RECT 51.800 96.800 52.200 97.200 ;
        RECT 54.200 96.800 54.600 97.200 ;
        RECT 55.000 96.800 55.400 97.200 ;
        RECT 59.800 96.800 60.200 97.200 ;
        RECT 30.200 95.800 30.600 96.200 ;
        RECT 33.400 95.800 33.800 96.200 ;
        RECT 27.000 94.800 27.400 95.200 ;
        RECT 29.400 94.800 29.800 95.200 ;
        RECT 22.200 93.800 22.600 94.200 ;
        RECT 24.600 93.800 25.000 94.200 ;
        RECT 26.200 93.800 26.600 94.200 ;
        RECT 24.600 93.200 24.900 93.800 ;
        RECT 27.000 93.200 27.300 94.800 ;
        RECT 11.800 92.800 12.200 93.200 ;
        RECT 12.600 92.800 13.000 93.200 ;
        RECT 20.600 92.800 21.000 93.200 ;
        RECT 24.600 92.800 25.000 93.200 ;
        RECT 25.400 92.800 25.800 93.200 ;
        RECT 27.000 92.800 27.400 93.200 ;
        RECT 25.400 92.200 25.700 92.800 ;
        RECT 25.400 91.800 25.800 92.200 ;
        RECT 25.400 90.800 25.800 91.200 ;
        RECT 14.200 89.800 14.600 90.200 ;
        RECT 14.200 89.200 14.500 89.800 ;
        RECT 25.400 89.200 25.700 90.800 ;
        RECT 14.200 88.800 14.600 89.200 ;
        RECT 15.800 88.800 16.200 89.200 ;
        RECT 21.400 89.100 21.800 89.200 ;
        RECT 22.200 89.100 22.600 89.200 ;
        RECT 21.400 88.800 22.600 89.100 ;
        RECT 25.400 88.800 25.800 89.200 ;
        RECT 11.800 87.100 12.200 87.200 ;
        RECT 12.600 87.100 13.000 87.200 ;
        RECT 11.800 86.800 13.000 87.100 ;
        RECT 12.600 85.800 13.000 86.200 ;
        RECT 14.200 86.100 14.600 86.200 ;
        RECT 15.000 86.100 15.400 86.200 ;
        RECT 14.200 85.800 15.400 86.100 ;
        RECT 12.600 82.200 12.900 85.800 ;
        RECT 15.800 85.200 16.100 88.800 ;
        RECT 20.700 87.800 21.100 87.900 ;
        RECT 20.700 87.500 23.500 87.800 ;
        RECT 23.800 87.500 24.200 87.900 ;
        RECT 17.400 86.800 17.800 87.200 ;
        RECT 18.200 86.800 18.600 87.200 ;
        RECT 19.800 86.800 20.200 87.200 ;
        RECT 17.400 86.200 17.700 86.800 ;
        RECT 18.200 86.200 18.500 86.800 ;
        RECT 17.400 85.800 17.800 86.200 ;
        RECT 18.200 85.800 18.600 86.200 ;
        RECT 15.000 85.100 15.400 85.200 ;
        RECT 15.800 85.100 16.200 85.200 ;
        RECT 15.000 84.800 16.200 85.100 ;
        RECT 16.600 84.800 17.000 85.200 ;
        RECT 15.800 83.800 16.200 84.200 ;
        RECT 12.600 81.800 13.000 82.200 ;
        RECT 15.800 79.200 16.100 83.800 ;
        RECT 16.600 82.200 16.900 84.800 ;
        RECT 16.600 81.800 17.000 82.200 ;
        RECT 17.400 81.200 17.700 85.800 ;
        RECT 19.800 85.200 20.100 86.800 ;
        RECT 19.800 84.800 20.200 85.200 ;
        RECT 20.700 85.100 21.000 87.500 ;
        RECT 21.400 87.400 21.800 87.500 ;
        RECT 23.100 87.400 23.500 87.500 ;
        RECT 23.900 87.100 24.200 87.500 ;
        RECT 21.400 86.800 24.200 87.100 ;
        RECT 24.600 87.100 25.000 87.200 ;
        RECT 25.400 87.100 25.800 87.200 ;
        RECT 24.600 86.800 25.800 87.100 ;
        RECT 27.000 86.800 27.400 87.200 ;
        RECT 21.400 86.100 21.700 86.800 ;
        RECT 21.300 85.700 21.700 86.100 ;
        RECT 23.900 85.100 24.200 86.800 ;
        RECT 27.000 86.200 27.300 86.800 ;
        RECT 20.700 84.700 21.100 85.100 ;
        RECT 23.800 84.700 24.200 85.100 ;
        RECT 25.400 85.800 25.800 86.200 ;
        RECT 27.000 85.800 27.400 86.200 ;
        RECT 27.800 85.800 28.200 86.200 ;
        RECT 28.600 85.800 29.000 86.200 ;
        RECT 25.400 85.200 25.700 85.800 ;
        RECT 25.400 84.800 25.800 85.200 ;
        RECT 18.200 84.100 18.600 84.200 ;
        RECT 19.000 84.100 19.400 84.200 ;
        RECT 18.200 83.800 19.400 84.100 ;
        RECT 17.400 80.800 17.800 81.200 ;
        RECT 27.000 79.200 27.300 85.800 ;
        RECT 27.800 85.200 28.100 85.800 ;
        RECT 28.600 85.200 28.900 85.800 ;
        RECT 29.400 85.200 29.700 94.800 ;
        RECT 30.200 93.200 30.500 95.800 ;
        RECT 31.800 95.100 32.200 95.200 ;
        RECT 32.600 95.100 33.000 95.200 ;
        RECT 31.800 94.800 33.000 95.100 ;
        RECT 30.200 92.800 30.600 93.200 ;
        RECT 33.400 92.200 33.700 95.800 ;
        RECT 34.200 93.200 34.500 96.800 ;
        RECT 37.400 95.800 37.800 96.200 ;
        RECT 42.200 96.100 42.600 96.200 ;
        RECT 40.600 95.800 42.600 96.100 ;
        RECT 45.400 95.800 45.800 96.200 ;
        RECT 35.000 94.800 35.400 95.200 ;
        RECT 35.800 94.800 36.200 95.200 ;
        RECT 36.600 94.800 37.000 95.200 ;
        RECT 35.000 94.200 35.300 94.800 ;
        RECT 35.800 94.200 36.100 94.800 ;
        RECT 36.600 94.200 36.900 94.800 ;
        RECT 37.400 94.200 37.700 95.800 ;
        RECT 38.200 95.100 38.600 95.200 ;
        RECT 39.000 95.100 39.400 95.200 ;
        RECT 38.200 94.800 39.400 95.100 ;
        RECT 40.600 94.200 40.900 95.800 ;
        RECT 43.000 94.800 43.400 95.200 ;
        RECT 35.000 93.800 35.400 94.200 ;
        RECT 35.800 93.800 36.200 94.200 ;
        RECT 36.600 93.800 37.000 94.200 ;
        RECT 37.400 93.800 37.800 94.200 ;
        RECT 40.600 93.800 41.000 94.200 ;
        RECT 41.400 94.100 41.800 94.200 ;
        RECT 42.200 94.100 42.600 94.200 ;
        RECT 41.400 93.800 42.600 94.100 ;
        RECT 34.200 92.800 34.600 93.200 ;
        RECT 33.400 92.100 33.800 92.200 ;
        RECT 32.600 91.800 33.800 92.100 ;
        RECT 30.200 87.800 30.600 88.200 ;
        RECT 30.200 87.200 30.500 87.800 ;
        RECT 30.200 86.800 30.600 87.200 ;
        RECT 32.600 86.200 32.900 91.800 ;
        RECT 41.400 89.200 41.700 93.800 ;
        RECT 37.400 89.100 37.800 89.200 ;
        RECT 36.600 88.800 37.800 89.100 ;
        RECT 41.400 88.800 41.800 89.200 ;
        RECT 33.400 87.100 33.800 87.200 ;
        RECT 34.200 87.100 34.600 87.200 ;
        RECT 33.400 86.800 34.600 87.100 ;
        RECT 30.200 85.800 30.600 86.200 ;
        RECT 32.600 85.800 33.000 86.200 ;
        RECT 34.200 85.800 34.600 86.200 ;
        RECT 35.800 85.800 36.200 86.200 ;
        RECT 27.800 84.800 28.200 85.200 ;
        RECT 28.600 84.800 29.000 85.200 ;
        RECT 29.400 84.800 29.800 85.200 ;
        RECT 14.200 78.800 14.600 79.200 ;
        RECT 15.800 78.800 16.200 79.200 ;
        RECT 27.000 78.800 27.400 79.200 ;
        RECT 12.600 76.100 13.000 76.200 ;
        RECT 13.400 76.100 13.800 76.200 ;
        RECT 12.600 75.800 13.800 76.100 ;
        RECT 12.600 75.200 12.900 75.800 ;
        RECT 14.200 75.200 14.500 78.800 ;
        RECT 15.000 76.800 15.400 77.200 ;
        RECT 19.800 76.800 20.200 77.200 ;
        RECT 12.600 74.800 13.000 75.200 ;
        RECT 14.200 74.800 14.600 75.200 ;
        RECT 11.800 73.800 12.200 74.200 ;
        RECT 11.800 73.200 12.100 73.800 ;
        RECT 11.800 72.800 12.200 73.200 ;
        RECT 12.600 69.200 12.900 74.800 ;
        RECT 15.000 74.200 15.300 76.800 ;
        RECT 19.800 76.200 20.100 76.800 ;
        RECT 16.600 76.100 17.000 76.200 ;
        RECT 17.400 76.100 17.800 76.200 ;
        RECT 16.600 75.800 17.800 76.100 ;
        RECT 19.800 75.800 20.200 76.200 ;
        RECT 21.400 75.800 21.800 76.200 ;
        RECT 24.600 76.100 25.000 76.200 ;
        RECT 25.400 76.100 25.800 76.200 ;
        RECT 24.600 75.800 25.800 76.100 ;
        RECT 27.000 76.100 27.400 76.200 ;
        RECT 27.800 76.100 28.200 76.200 ;
        RECT 27.000 75.800 28.200 76.100 ;
        RECT 19.800 75.100 20.200 75.200 ;
        RECT 20.600 75.100 21.000 75.200 ;
        RECT 19.800 74.800 21.000 75.100 ;
        RECT 13.400 73.800 13.800 74.200 ;
        RECT 15.000 73.800 15.400 74.200 ;
        RECT 18.200 73.800 18.600 74.200 ;
        RECT 19.000 73.800 19.400 74.200 ;
        RECT 11.000 68.800 11.400 69.200 ;
        RECT 12.600 68.800 13.000 69.200 ;
        RECT 3.000 67.800 3.400 68.200 ;
        RECT 4.600 67.800 5.000 68.200 ;
        RECT 5.400 67.800 5.800 68.200 ;
        RECT 5.400 66.200 5.700 67.800 ;
        RECT 7.800 67.100 8.200 67.200 ;
        RECT 8.600 67.100 9.000 67.200 ;
        RECT 7.800 66.800 9.000 67.100 ;
        RECT 11.000 66.800 11.400 67.200 ;
        RECT 5.400 65.800 5.800 66.200 ;
        RECT 8.600 65.800 9.000 66.200 ;
        RECT 9.400 65.800 9.800 66.200 ;
        RECT 10.200 65.800 10.600 66.200 ;
        RECT 8.600 65.200 8.900 65.800 ;
        RECT 9.400 65.200 9.700 65.800 ;
        RECT 10.200 65.200 10.500 65.800 ;
        RECT 2.200 64.800 2.600 65.200 ;
        RECT 6.200 64.800 6.600 65.200 ;
        RECT 8.600 64.800 9.000 65.200 ;
        RECT 9.400 64.800 9.800 65.200 ;
        RECT 10.200 64.800 10.600 65.200 ;
        RECT 5.400 57.800 5.800 58.200 ;
        RECT 5.400 57.200 5.700 57.800 ;
        RECT 3.800 57.100 4.200 57.200 ;
        RECT 4.600 57.100 5.000 57.200 ;
        RECT 3.800 56.800 5.000 57.100 ;
        RECT 5.400 56.800 5.800 57.200 ;
        RECT 3.000 55.100 3.400 55.200 ;
        RECT 3.800 55.100 4.200 55.200 ;
        RECT 3.000 54.800 4.200 55.100 ;
        RECT 3.800 51.800 4.200 52.200 ;
        RECT 2.200 47.800 2.600 48.200 ;
        RECT 2.200 47.000 2.500 47.800 ;
        RECT 3.800 47.200 4.100 51.800 ;
        RECT 6.200 49.200 6.500 64.800 ;
        RECT 8.600 63.800 9.000 64.200 ;
        RECT 7.800 62.800 8.200 63.200 ;
        RECT 7.000 53.800 7.400 54.200 ;
        RECT 7.000 49.200 7.300 53.800 ;
        RECT 7.800 53.200 8.100 62.800 ;
        RECT 8.600 57.200 8.900 63.800 ;
        RECT 10.200 57.200 10.500 64.800 ;
        RECT 11.000 64.200 11.300 66.800 ;
        RECT 11.800 64.800 12.200 65.200 ;
        RECT 11.000 63.800 11.400 64.200 ;
        RECT 8.600 56.800 9.000 57.200 ;
        RECT 10.200 56.800 10.600 57.200 ;
        RECT 11.000 56.100 11.300 63.800 ;
        RECT 11.800 57.200 12.100 64.800 ;
        RECT 13.400 59.200 13.700 73.800 ;
        RECT 18.200 73.200 18.500 73.800 ;
        RECT 16.600 72.800 17.000 73.200 ;
        RECT 17.400 72.800 17.800 73.200 ;
        RECT 18.200 72.800 18.600 73.200 ;
        RECT 15.000 70.800 15.400 71.200 ;
        RECT 14.200 65.800 14.600 66.200 ;
        RECT 14.200 64.200 14.500 65.800 ;
        RECT 15.000 65.200 15.300 70.800 ;
        RECT 16.600 69.200 16.900 72.800 ;
        RECT 16.600 68.800 17.000 69.200 ;
        RECT 15.800 66.100 16.200 66.200 ;
        RECT 16.600 66.100 17.000 66.200 ;
        RECT 15.800 65.800 17.000 66.100 ;
        RECT 17.400 65.200 17.700 72.800 ;
        RECT 19.000 66.200 19.300 73.800 ;
        RECT 21.400 72.200 21.700 75.800 ;
        RECT 23.000 74.800 23.400 75.200 ;
        RECT 27.000 74.800 27.400 75.200 ;
        RECT 29.400 74.800 29.800 75.200 ;
        RECT 22.200 73.800 22.600 74.200 ;
        RECT 22.200 73.200 22.500 73.800 ;
        RECT 22.200 72.800 22.600 73.200 ;
        RECT 21.400 71.800 21.800 72.200 ;
        RECT 23.000 69.200 23.300 74.800 ;
        RECT 27.000 74.200 27.300 74.800 ;
        RECT 29.400 74.200 29.700 74.800 ;
        RECT 27.000 73.800 27.400 74.200 ;
        RECT 29.400 73.800 29.800 74.200 ;
        RECT 25.400 72.800 25.800 73.200 ;
        RECT 26.200 72.800 26.600 73.200 ;
        RECT 27.000 73.100 27.400 73.200 ;
        RECT 27.800 73.100 28.200 73.200 ;
        RECT 27.000 72.800 28.200 73.100 ;
        RECT 25.400 72.200 25.700 72.800 ;
        RECT 25.400 71.800 25.800 72.200 ;
        RECT 20.600 68.800 21.000 69.200 ;
        RECT 22.200 68.800 22.600 69.200 ;
        RECT 23.000 68.800 23.400 69.200 ;
        RECT 20.600 66.200 20.900 68.800 ;
        RECT 21.400 67.800 21.800 68.200 ;
        RECT 21.400 67.200 21.700 67.800 ;
        RECT 21.400 66.800 21.800 67.200 ;
        RECT 22.200 66.200 22.500 68.800 ;
        RECT 23.800 68.100 24.200 68.200 ;
        RECT 24.600 68.100 25.000 68.200 ;
        RECT 23.800 67.800 25.000 68.100 ;
        RECT 23.800 66.800 24.200 67.200 ;
        RECT 23.800 66.200 24.100 66.800 ;
        RECT 25.400 66.200 25.700 71.800 ;
        RECT 26.200 71.200 26.500 72.800 ;
        RECT 26.200 70.800 26.600 71.200 ;
        RECT 27.800 69.800 28.200 70.200 ;
        RECT 27.800 67.200 28.100 69.800 ;
        RECT 30.200 69.200 30.500 85.800 ;
        RECT 34.200 85.200 34.500 85.800 ;
        RECT 35.800 85.200 36.100 85.800 ;
        RECT 36.600 85.200 36.900 88.800 ;
        RECT 37.400 88.200 37.700 88.800 ;
        RECT 37.400 87.800 37.800 88.200 ;
        RECT 40.600 87.800 41.000 88.200 ;
        RECT 40.600 87.200 40.900 87.800 ;
        RECT 43.000 87.200 43.300 94.800 ;
        RECT 45.400 92.200 45.700 95.800 ;
        RECT 46.200 95.200 46.500 96.800 ;
        RECT 50.200 95.800 50.600 96.200 ;
        RECT 46.200 94.800 46.600 95.200 ;
        RECT 50.200 94.100 50.500 95.800 ;
        RECT 51.000 95.200 51.300 96.800 ;
        RECT 53.400 95.800 53.800 96.200 ;
        RECT 54.200 95.800 54.600 96.200 ;
        RECT 51.000 94.800 51.400 95.200 ;
        RECT 53.400 94.200 53.700 95.800 ;
        RECT 54.200 95.200 54.500 95.800 ;
        RECT 54.200 94.800 54.600 95.200 ;
        RECT 50.200 93.800 51.300 94.100 ;
        RECT 53.400 93.800 53.800 94.200 ;
        RECT 50.200 93.200 50.500 93.800 ;
        RECT 50.200 92.800 50.600 93.200 ;
        RECT 43.800 91.800 44.200 92.200 ;
        RECT 45.400 91.800 45.800 92.200 ;
        RECT 43.800 89.200 44.100 91.800 ;
        RECT 51.000 89.200 51.300 93.800 ;
        RECT 55.000 92.200 55.300 96.800 ;
        RECT 56.600 94.800 57.000 95.200 ;
        RECT 55.000 91.800 55.400 92.200 ;
        RECT 43.800 88.800 44.200 89.200 ;
        RECT 44.600 88.800 45.000 89.200 ;
        RECT 51.000 88.800 51.400 89.200 ;
        RECT 54.200 88.800 54.600 89.200 ;
        RECT 44.600 87.200 44.900 88.800 ;
        RECT 37.400 87.100 37.800 87.200 ;
        RECT 38.200 87.100 38.600 87.200 ;
        RECT 37.400 86.800 38.600 87.100 ;
        RECT 39.000 87.100 39.400 87.200 ;
        RECT 39.800 87.100 40.200 87.200 ;
        RECT 39.000 86.800 40.200 87.100 ;
        RECT 40.600 86.800 41.000 87.200 ;
        RECT 43.000 86.800 43.400 87.200 ;
        RECT 44.600 86.800 45.000 87.200 ;
        RECT 47.800 87.100 48.200 87.200 ;
        RECT 48.600 87.100 49.000 87.200 ;
        RECT 47.800 86.800 49.000 87.100 ;
        RECT 50.200 86.800 50.600 87.200 ;
        RECT 52.600 87.100 53.000 87.200 ;
        RECT 53.400 87.100 53.800 87.200 ;
        RECT 52.600 86.800 53.800 87.100 ;
        RECT 39.000 86.100 39.400 86.200 ;
        RECT 39.800 86.100 40.200 86.200 ;
        RECT 39.000 85.800 40.200 86.100 ;
        RECT 44.600 85.800 45.000 86.200 ;
        RECT 47.800 85.800 48.200 86.200 ;
        RECT 44.600 85.200 44.900 85.800 ;
        RECT 47.800 85.200 48.100 85.800 ;
        RECT 31.000 85.100 31.400 85.200 ;
        RECT 31.800 85.100 32.200 85.200 ;
        RECT 31.000 84.800 32.200 85.100 ;
        RECT 34.200 84.800 34.600 85.200 ;
        RECT 35.800 84.800 36.200 85.200 ;
        RECT 36.600 84.800 37.000 85.200 ;
        RECT 43.000 85.100 43.400 85.200 ;
        RECT 43.800 85.100 44.200 85.200 ;
        RECT 43.000 84.800 44.200 85.100 ;
        RECT 44.600 84.800 45.000 85.200 ;
        RECT 45.400 84.800 45.800 85.200 ;
        RECT 47.800 84.800 48.200 85.200 ;
        RECT 32.600 83.800 33.000 84.200 ;
        RECT 35.000 84.100 35.400 84.200 ;
        RECT 35.800 84.100 36.200 84.200 ;
        RECT 35.000 83.800 36.200 84.100 ;
        RECT 32.600 83.200 32.900 83.800 ;
        RECT 32.600 82.800 33.000 83.200 ;
        RECT 45.400 78.200 45.700 84.800 ;
        RECT 50.200 79.200 50.500 86.800 ;
        RECT 52.600 85.800 53.000 86.200 ;
        RECT 52.600 85.200 52.900 85.800 ;
        RECT 51.800 84.800 52.200 85.200 ;
        RECT 52.600 84.800 53.000 85.200 ;
        RECT 53.400 84.800 53.800 85.200 ;
        RECT 51.800 84.200 52.100 84.800 ;
        RECT 53.400 84.200 53.700 84.800 ;
        RECT 51.800 83.800 52.200 84.200 ;
        RECT 53.400 83.800 53.800 84.200 ;
        RECT 53.400 80.800 53.800 81.200 ;
        RECT 51.000 79.800 51.400 80.200 ;
        RECT 50.200 78.800 50.600 79.200 ;
        RECT 43.000 77.800 43.400 78.200 ;
        RECT 45.400 77.800 45.800 78.200 ;
        RECT 49.400 77.800 49.800 78.200 ;
        RECT 43.000 77.200 43.300 77.800 ;
        RECT 33.400 76.800 33.800 77.200 ;
        RECT 42.200 76.800 42.600 77.200 ;
        RECT 43.000 76.800 43.400 77.200 ;
        RECT 33.400 76.200 33.700 76.800 ;
        RECT 33.400 75.800 33.800 76.200 ;
        RECT 35.000 75.800 35.400 76.200 ;
        RECT 33.400 74.800 33.800 75.200 ;
        RECT 33.400 74.200 33.700 74.800 ;
        RECT 31.800 73.800 32.200 74.200 ;
        RECT 33.400 73.800 33.800 74.200 ;
        RECT 31.800 69.200 32.100 73.800 ;
        RECT 34.200 72.800 34.600 73.200 ;
        RECT 34.200 70.200 34.500 72.800 ;
        RECT 35.000 72.200 35.300 75.800 ;
        RECT 38.200 74.100 38.600 74.200 ;
        RECT 39.000 74.100 39.400 74.200 ;
        RECT 38.200 73.800 39.400 74.100 ;
        RECT 42.200 73.200 42.500 76.800 ;
        RECT 49.400 76.200 49.700 77.800 ;
        RECT 51.000 77.200 51.300 79.800 ;
        RECT 52.600 77.800 53.000 78.200 ;
        RECT 52.600 77.200 52.900 77.800 ;
        RECT 50.200 76.800 50.600 77.200 ;
        RECT 51.000 76.800 51.400 77.200 ;
        RECT 52.600 76.800 53.000 77.200 ;
        RECT 49.400 75.800 49.800 76.200 ;
        RECT 50.200 75.200 50.500 76.800 ;
        RECT 53.400 76.200 53.700 80.800 ;
        RECT 54.200 80.100 54.500 88.800 ;
        RECT 56.600 88.200 56.900 94.800 ;
        RECT 59.800 94.200 60.100 96.800 ;
        RECT 61.400 95.800 61.800 96.200 ;
        RECT 60.600 94.800 61.000 95.200 ;
        RECT 61.400 95.100 61.700 95.800 ;
        RECT 62.200 95.100 62.600 95.200 ;
        RECT 61.400 94.800 62.600 95.100 ;
        RECT 59.800 93.800 60.200 94.200 ;
        RECT 58.200 93.100 58.600 93.200 ;
        RECT 58.200 92.800 59.300 93.100 ;
        RECT 59.000 89.200 59.300 92.800 ;
        RECT 59.000 88.800 59.400 89.200 ;
        RECT 56.600 87.800 57.000 88.200 ;
        RECT 57.400 87.800 57.800 88.200 ;
        RECT 58.200 88.100 58.600 88.200 ;
        RECT 59.000 88.100 59.400 88.200 ;
        RECT 58.200 87.800 59.400 88.100 ;
        RECT 57.400 87.200 57.700 87.800 ;
        RECT 57.400 86.800 57.800 87.200 ;
        RECT 55.000 84.800 55.400 85.200 ;
        RECT 55.000 81.200 55.300 84.800 ;
        RECT 55.000 80.800 55.400 81.200 ;
        RECT 54.200 79.800 55.300 80.100 ;
        RECT 55.000 79.200 55.300 79.800 ;
        RECT 55.800 79.800 56.200 80.200 ;
        RECT 55.000 78.800 55.400 79.200 ;
        RECT 55.800 78.200 56.100 79.800 ;
        RECT 58.200 79.100 58.500 87.800 ;
        RECT 59.800 84.200 60.100 93.800 ;
        RECT 60.600 92.200 60.900 94.800 ;
        RECT 62.200 93.200 62.500 94.800 ;
        RECT 62.200 92.800 62.600 93.200 ;
        RECT 60.600 91.800 61.000 92.200 ;
        RECT 63.000 89.200 63.300 105.800 ;
        RECT 63.800 105.200 64.100 105.800 ;
        RECT 67.000 105.200 67.300 114.800 ;
        RECT 67.800 113.800 68.200 114.200 ;
        RECT 67.800 107.200 68.100 113.800 ;
        RECT 69.400 113.200 69.700 116.800 ;
        RECT 73.400 115.800 73.800 116.200 ;
        RECT 76.600 115.800 77.000 116.200 ;
        RECT 70.200 115.100 70.600 115.200 ;
        RECT 71.000 115.100 71.400 115.200 ;
        RECT 70.200 114.800 71.400 115.100 ;
        RECT 71.800 114.800 72.200 115.200 ;
        RECT 71.000 113.800 71.400 114.200 ;
        RECT 69.400 112.800 69.800 113.200 ;
        RECT 71.000 112.200 71.300 113.800 ;
        RECT 71.000 111.800 71.400 112.200 ;
        RECT 71.000 107.800 71.400 108.200 ;
        RECT 67.800 106.800 68.200 107.200 ;
        RECT 68.600 107.100 69.000 107.200 ;
        RECT 69.400 107.100 69.800 107.200 ;
        RECT 68.600 106.800 69.800 107.100 ;
        RECT 67.800 106.200 68.100 106.800 ;
        RECT 71.000 106.200 71.300 107.800 ;
        RECT 71.800 107.200 72.100 114.800 ;
        RECT 73.400 114.200 73.700 115.800 ;
        RECT 75.000 115.100 75.400 115.200 ;
        RECT 75.800 115.100 76.200 115.200 ;
        RECT 75.000 114.800 76.200 115.100 ;
        RECT 73.400 113.800 73.800 114.200 ;
        RECT 76.600 109.200 76.900 115.800 ;
        RECT 79.000 115.200 79.300 119.800 ;
        RECT 80.600 115.200 80.900 123.800 ;
        RECT 81.400 121.800 81.800 122.200 ;
        RECT 81.400 118.200 81.700 121.800 ;
        RECT 81.400 117.800 81.800 118.200 ;
        RECT 81.400 115.800 81.800 116.200 ;
        RECT 77.400 114.800 77.800 115.200 ;
        RECT 79.000 114.800 79.400 115.200 ;
        RECT 80.600 114.800 81.000 115.200 ;
        RECT 77.400 113.200 77.700 114.800 ;
        RECT 77.400 112.800 77.800 113.200 ;
        RECT 80.600 111.800 81.000 112.200 ;
        RECT 80.600 109.200 80.900 111.800 ;
        RECT 81.400 111.200 81.700 115.800 ;
        RECT 84.600 115.200 84.900 125.800 ;
        RECT 87.000 122.100 87.400 128.900 ;
        RECT 87.800 122.100 88.200 128.900 ;
        RECT 88.600 123.100 89.000 128.900 ;
        RECT 89.400 126.800 89.800 127.200 ;
        RECT 89.400 126.200 89.700 126.800 ;
        RECT 89.400 125.800 89.800 126.200 ;
        RECT 90.200 123.100 90.600 128.900 ;
        RECT 91.800 123.100 92.200 128.900 ;
        RECT 92.600 122.100 93.000 128.900 ;
        RECT 93.400 122.100 93.800 128.900 ;
        RECT 94.200 122.100 94.600 128.900 ;
        RECT 95.000 126.800 95.400 127.200 ;
        RECT 95.000 126.200 95.300 126.800 ;
        RECT 95.000 125.800 95.400 126.200 ;
        RECT 103.000 126.100 103.400 126.200 ;
        RECT 103.800 126.100 104.200 126.200 ;
        RECT 103.000 125.800 104.200 126.100 ;
        RECT 103.000 124.800 103.400 125.200 ;
        RECT 99.000 122.100 99.400 122.200 ;
        RECT 99.800 122.100 100.200 122.200 ;
        RECT 99.000 121.800 100.200 122.100 ;
        RECT 84.600 114.800 85.000 115.200 ;
        RECT 83.800 112.800 84.200 113.200 ;
        RECT 81.400 110.800 81.800 111.200 ;
        RECT 83.800 109.200 84.100 112.800 ;
        RECT 86.200 112.100 86.600 118.900 ;
        RECT 87.000 112.100 87.400 118.900 ;
        RECT 87.800 112.100 88.200 117.900 ;
        RECT 88.600 113.800 89.000 114.200 ;
        RECT 87.000 110.800 87.400 111.200 ;
        RECT 88.600 111.100 88.900 113.800 ;
        RECT 89.400 112.100 89.800 117.900 ;
        RECT 91.000 112.100 91.400 117.900 ;
        RECT 91.800 112.100 92.200 118.900 ;
        RECT 92.600 112.100 93.000 118.900 ;
        RECT 93.400 112.100 93.800 118.900 ;
        RECT 99.800 115.200 100.100 121.800 ;
        RECT 101.400 117.100 101.800 117.200 ;
        RECT 102.200 117.100 102.600 117.200 ;
        RECT 101.400 116.800 102.600 117.100 ;
        RECT 99.800 114.800 100.200 115.200 ;
        RECT 98.200 112.800 98.600 113.200 ;
        RECT 98.200 112.200 98.500 112.800 ;
        RECT 99.800 112.200 100.100 114.800 ;
        RECT 103.000 113.200 103.300 124.800 ;
        RECT 106.200 122.100 106.600 128.900 ;
        RECT 107.000 122.100 107.400 128.900 ;
        RECT 107.800 123.100 108.200 128.900 ;
        RECT 108.600 126.800 109.000 127.200 ;
        RECT 108.600 119.200 108.900 126.800 ;
        RECT 109.400 123.100 109.800 128.900 ;
        RECT 111.000 123.100 111.400 128.900 ;
        RECT 111.800 122.100 112.200 128.900 ;
        RECT 112.600 122.100 113.000 128.900 ;
        RECT 113.400 122.100 113.800 128.900 ;
        RECT 120.600 128.100 121.000 128.200 ;
        RECT 121.400 128.100 121.800 128.200 ;
        RECT 120.600 127.800 121.800 128.100 ;
        RECT 122.200 126.100 122.600 126.200 ;
        RECT 123.000 126.100 123.400 126.200 ;
        RECT 122.200 125.800 123.400 126.100 ;
        RECT 124.600 125.800 125.000 126.200 ;
        RECT 118.200 121.800 118.600 122.200 ;
        RECT 119.800 121.800 120.200 122.200 ;
        RECT 118.200 121.200 118.500 121.800 ;
        RECT 113.400 120.800 113.800 121.200 ;
        RECT 118.200 120.800 118.600 121.200 ;
        RECT 105.400 118.800 105.800 119.200 ;
        RECT 106.200 119.100 106.600 119.200 ;
        RECT 107.000 119.100 107.400 119.200 ;
        RECT 106.200 118.800 107.400 119.100 ;
        RECT 108.600 118.800 109.000 119.200 ;
        RECT 105.400 116.100 105.700 118.800 ;
        RECT 109.400 117.100 109.800 117.200 ;
        RECT 110.200 117.100 110.600 117.200 ;
        RECT 109.400 116.800 110.600 117.100 ;
        RECT 111.000 116.800 111.400 117.200 ;
        RECT 111.000 116.200 111.300 116.800 ;
        RECT 105.400 115.800 106.500 116.100 ;
        RECT 104.600 115.100 105.000 115.200 ;
        RECT 105.400 115.100 105.800 115.200 ;
        RECT 104.600 114.800 105.800 115.100 ;
        RECT 106.200 114.200 106.500 115.800 ;
        RECT 108.600 115.800 109.000 116.200 ;
        RECT 111.000 115.800 111.400 116.200 ;
        RECT 111.800 116.100 112.200 116.200 ;
        RECT 112.600 116.100 113.000 116.200 ;
        RECT 111.800 115.800 113.000 116.100 ;
        RECT 108.600 115.200 108.900 115.800 ;
        RECT 111.000 115.200 111.300 115.800 ;
        RECT 108.600 114.800 109.000 115.200 ;
        RECT 111.000 114.800 111.400 115.200 ;
        RECT 104.600 114.100 105.000 114.200 ;
        RECT 105.400 114.100 105.800 114.200 ;
        RECT 104.600 113.800 105.800 114.100 ;
        RECT 106.200 113.800 106.600 114.200 ;
        RECT 107.000 114.100 107.400 114.200 ;
        RECT 107.800 114.100 108.200 114.200 ;
        RECT 107.000 113.800 108.200 114.100 ;
        RECT 113.400 113.200 113.700 120.800 ;
        RECT 116.600 119.800 117.000 120.200 ;
        RECT 116.600 119.200 116.900 119.800 ;
        RECT 116.600 118.800 117.000 119.200 ;
        RECT 119.800 116.200 120.100 121.800 ;
        RECT 114.200 115.800 114.600 116.200 ;
        RECT 119.800 115.800 120.200 116.200 ;
        RECT 120.600 116.100 121.000 116.200 ;
        RECT 121.400 116.100 121.800 116.200 ;
        RECT 120.600 115.800 121.800 116.100 ;
        RECT 114.200 115.200 114.500 115.800 ;
        RECT 124.600 115.200 124.900 125.800 ;
        RECT 125.400 122.100 125.800 128.900 ;
        RECT 126.200 122.100 126.600 128.900 ;
        RECT 127.000 123.100 127.400 128.900 ;
        RECT 127.800 126.800 128.200 127.200 ;
        RECT 127.800 120.200 128.100 126.800 ;
        RECT 128.600 123.100 129.000 128.900 ;
        RECT 130.200 123.100 130.600 128.900 ;
        RECT 131.000 122.100 131.400 128.900 ;
        RECT 131.800 122.100 132.200 128.900 ;
        RECT 132.600 122.100 133.000 128.900 ;
        RECT 137.400 128.100 137.800 128.200 ;
        RECT 138.200 128.100 138.600 128.200 ;
        RECT 137.400 127.800 138.600 128.100 ;
        RECT 141.400 125.800 141.800 126.200 ;
        RECT 143.800 125.800 144.200 126.200 ;
        RECT 141.400 122.200 141.700 125.800 ;
        RECT 143.800 125.200 144.100 125.800 ;
        RECT 143.800 124.800 144.200 125.200 ;
        RECT 147.800 124.800 148.200 125.200 ;
        RECT 147.800 124.200 148.100 124.800 ;
        RECT 147.800 123.800 148.200 124.200 ;
        RECT 141.400 121.800 141.800 122.200 ;
        RECT 147.000 121.800 147.400 122.200 ;
        RECT 148.600 121.800 149.000 122.200 ;
        RECT 140.600 120.800 141.000 121.200 ;
        RECT 127.800 119.800 128.200 120.200 ;
        RECT 114.200 114.800 114.600 115.200 ;
        RECT 116.600 114.800 117.000 115.200 ;
        RECT 117.400 114.800 117.800 115.200 ;
        RECT 118.200 114.800 118.600 115.200 ;
        RECT 120.600 114.800 121.000 115.200 ;
        RECT 121.400 115.100 121.800 115.200 ;
        RECT 121.400 114.800 122.500 115.100 ;
        RECT 116.600 114.200 116.900 114.800 ;
        RECT 117.400 114.200 117.700 114.800 ;
        RECT 114.200 114.100 114.600 114.200 ;
        RECT 115.000 114.100 115.400 114.200 ;
        RECT 114.200 113.800 115.400 114.100 ;
        RECT 116.600 113.800 117.000 114.200 ;
        RECT 117.400 113.800 117.800 114.200 ;
        RECT 118.200 113.200 118.500 114.800 ;
        RECT 120.600 114.200 120.900 114.800 ;
        RECT 119.000 114.100 119.400 114.200 ;
        RECT 119.800 114.100 120.200 114.200 ;
        RECT 119.000 113.800 120.200 114.100 ;
        RECT 120.600 113.800 121.000 114.200 ;
        RECT 102.200 113.100 102.600 113.200 ;
        RECT 103.000 113.100 103.400 113.200 ;
        RECT 102.200 112.800 103.400 113.100 ;
        RECT 113.400 112.800 113.800 113.200 ;
        RECT 118.200 112.800 118.600 113.200 ;
        RECT 95.800 111.800 96.200 112.200 ;
        RECT 98.200 111.800 98.600 112.200 ;
        RECT 99.800 111.800 100.200 112.200 ;
        RECT 111.000 111.800 111.400 112.200 ;
        RECT 88.600 110.800 89.700 111.100 ;
        RECT 87.000 109.200 87.300 110.800 ;
        RECT 89.400 109.200 89.700 110.800 ;
        RECT 92.600 110.800 93.000 111.200 ;
        RECT 91.800 109.800 92.200 110.200 ;
        RECT 76.600 108.800 77.000 109.200 ;
        RECT 80.600 108.800 81.000 109.200 ;
        RECT 83.800 108.800 84.200 109.200 ;
        RECT 86.200 108.800 86.600 109.200 ;
        RECT 87.000 108.800 87.400 109.200 ;
        RECT 89.400 108.800 89.800 109.200 ;
        RECT 86.200 108.200 86.500 108.800 ;
        RECT 72.600 108.100 73.000 108.200 ;
        RECT 73.400 108.100 73.800 108.200 ;
        RECT 72.600 107.800 73.800 108.100 ;
        RECT 78.200 107.800 78.600 108.200 ;
        RECT 79.800 107.800 80.200 108.200 ;
        RECT 86.200 107.800 86.600 108.200 ;
        RECT 90.200 108.100 90.600 108.200 ;
        RECT 91.000 108.100 91.400 108.200 ;
        RECT 90.200 107.800 91.400 108.100 ;
        RECT 78.200 107.200 78.500 107.800 ;
        RECT 71.800 106.800 72.200 107.200 ;
        RECT 72.600 107.100 73.000 107.200 ;
        RECT 73.400 107.100 73.800 107.200 ;
        RECT 72.600 106.800 73.800 107.100 ;
        RECT 74.200 106.800 74.600 107.200 ;
        RECT 75.800 107.100 76.200 107.200 ;
        RECT 75.800 106.800 76.900 107.100 ;
        RECT 78.200 106.800 78.600 107.200 ;
        RECT 74.200 106.200 74.500 106.800 ;
        RECT 67.800 105.800 68.200 106.200 ;
        RECT 69.400 105.800 69.800 106.200 ;
        RECT 70.200 105.800 70.600 106.200 ;
        RECT 71.000 105.800 71.400 106.200 ;
        RECT 74.200 105.800 74.600 106.200 ;
        RECT 75.000 105.800 75.400 106.200 ;
        RECT 75.800 105.800 76.200 106.200 ;
        RECT 69.400 105.200 69.700 105.800 ;
        RECT 63.800 104.800 64.200 105.200 ;
        RECT 64.600 105.100 65.000 105.200 ;
        RECT 65.400 105.100 65.800 105.200 ;
        RECT 64.600 104.800 65.800 105.100 ;
        RECT 66.200 105.100 66.600 105.200 ;
        RECT 67.000 105.100 67.400 105.200 ;
        RECT 66.200 104.800 67.400 105.100 ;
        RECT 69.400 104.800 69.800 105.200 ;
        RECT 70.200 104.200 70.500 105.800 ;
        RECT 75.000 105.200 75.300 105.800 ;
        RECT 75.800 105.200 76.100 105.800 ;
        RECT 71.800 105.100 72.200 105.200 ;
        RECT 72.600 105.100 73.000 105.200 ;
        RECT 71.800 104.800 73.000 105.100 ;
        RECT 75.000 104.800 75.400 105.200 ;
        RECT 75.800 104.800 76.200 105.200 ;
        RECT 70.200 103.800 70.600 104.200 ;
        RECT 69.400 102.800 69.800 103.200 ;
        RECT 65.400 101.800 65.800 102.200 ;
        RECT 65.400 99.200 65.700 101.800 ;
        RECT 69.400 99.200 69.700 102.800 ;
        RECT 65.400 98.800 65.800 99.200 ;
        RECT 69.400 98.800 69.800 99.200 ;
        RECT 65.400 96.800 65.800 97.200 ;
        RECT 70.200 97.100 70.600 97.200 ;
        RECT 71.000 97.100 71.400 97.200 ;
        RECT 70.200 96.800 71.400 97.100 ;
        RECT 64.600 94.800 65.000 95.200 ;
        RECT 64.600 94.200 64.900 94.800 ;
        RECT 63.800 93.800 64.200 94.200 ;
        RECT 64.600 93.800 65.000 94.200 ;
        RECT 63.800 93.200 64.100 93.800 ;
        RECT 63.800 92.800 64.200 93.200 ;
        RECT 64.600 92.200 64.900 93.800 ;
        RECT 65.400 93.200 65.700 96.800 ;
        RECT 76.600 96.200 76.900 106.800 ;
        RECT 77.400 104.800 77.800 105.200 ;
        RECT 77.400 98.200 77.700 104.800 ;
        RECT 79.800 102.200 80.100 107.800 ;
        RECT 91.800 107.200 92.100 109.800 ;
        RECT 92.600 109.200 92.900 110.800 ;
        RECT 92.600 108.800 93.000 109.200 ;
        RECT 95.800 108.200 96.100 111.800 ;
        RECT 98.200 108.200 98.500 111.800 ;
        RECT 111.000 110.200 111.300 111.800 ;
        RECT 111.000 109.800 111.400 110.200 ;
        RECT 99.800 108.800 100.200 109.200 ;
        RECT 99.800 108.200 100.100 108.800 ;
        RECT 95.800 107.800 96.200 108.200 ;
        RECT 96.600 107.800 97.000 108.200 ;
        RECT 98.200 107.800 98.600 108.200 ;
        RECT 99.000 107.800 99.400 108.200 ;
        RECT 99.800 107.800 100.200 108.200 ;
        RECT 96.600 107.200 96.900 107.800 ;
        RECT 81.400 106.800 81.800 107.200 ;
        RECT 87.800 107.100 88.200 107.200 ;
        RECT 88.600 107.100 89.000 107.200 ;
        RECT 87.800 106.800 89.000 107.100 ;
        RECT 91.800 106.800 92.200 107.200 ;
        RECT 96.600 106.800 97.000 107.200 ;
        RECT 81.400 104.200 81.700 106.800 ;
        RECT 82.200 105.800 82.600 106.200 ;
        RECT 83.000 106.100 83.400 106.200 ;
        RECT 83.800 106.100 84.200 106.200 ;
        RECT 83.000 105.800 84.200 106.100 ;
        RECT 87.800 105.800 88.200 106.200 ;
        RECT 91.000 106.100 91.400 106.200 ;
        RECT 91.800 106.100 92.200 106.200 ;
        RECT 91.000 105.800 92.200 106.100 ;
        RECT 81.400 103.800 81.800 104.200 ;
        RECT 79.800 101.800 80.200 102.200 ;
        RECT 82.200 99.200 82.500 105.800 ;
        RECT 83.000 104.800 83.400 105.200 ;
        RECT 83.800 104.800 84.200 105.200 ;
        RECT 83.000 99.200 83.300 104.800 ;
        RECT 83.800 102.200 84.100 104.800 ;
        RECT 84.600 104.100 85.000 104.200 ;
        RECT 85.400 104.100 85.800 104.200 ;
        RECT 84.600 103.800 85.800 104.100 ;
        RECT 87.800 103.200 88.100 105.800 ;
        RECT 91.000 103.800 91.400 104.200 ;
        RECT 87.800 102.800 88.200 103.200 ;
        RECT 83.800 101.800 84.200 102.200 ;
        RECT 87.000 101.800 87.400 102.200 ;
        RECT 87.800 101.800 88.200 102.200 ;
        RECT 82.200 98.800 82.600 99.200 ;
        RECT 83.000 98.800 83.400 99.200 ;
        RECT 85.400 99.100 85.800 99.200 ;
        RECT 86.200 99.100 86.600 99.200 ;
        RECT 85.400 98.800 86.600 99.100 ;
        RECT 77.400 97.800 77.800 98.200 ;
        RECT 67.800 95.800 68.200 96.200 ;
        RECT 68.600 95.800 69.000 96.200 ;
        RECT 69.400 95.800 69.800 96.200 ;
        RECT 74.200 95.800 74.600 96.200 ;
        RECT 76.600 95.800 77.000 96.200 ;
        RECT 67.800 95.200 68.100 95.800 ;
        RECT 67.800 94.800 68.200 95.200 ;
        RECT 67.000 93.800 67.400 94.200 ;
        RECT 67.800 94.100 68.200 94.200 ;
        RECT 68.600 94.100 68.900 95.800 ;
        RECT 67.800 93.800 68.900 94.100 ;
        RECT 65.400 92.800 65.800 93.200 ;
        RECT 64.600 91.800 65.000 92.200 ;
        RECT 63.800 90.800 64.200 91.200 ;
        RECT 63.800 89.200 64.100 90.800 ;
        RECT 67.000 89.200 67.300 93.800 ;
        RECT 63.000 88.800 63.400 89.200 ;
        RECT 63.800 88.800 64.200 89.200 ;
        RECT 67.000 88.800 67.400 89.200 ;
        RECT 61.400 87.800 61.800 88.200 ;
        RECT 61.400 87.200 61.700 87.800 ;
        RECT 61.400 86.800 61.800 87.200 ;
        RECT 66.200 86.800 66.600 87.200 ;
        RECT 63.800 85.800 64.200 86.200 ;
        RECT 65.400 85.800 65.800 86.200 ;
        RECT 63.800 85.200 64.100 85.800 ;
        RECT 63.800 84.800 64.200 85.200 ;
        RECT 59.800 83.800 60.200 84.200 ;
        RECT 64.600 83.800 65.000 84.200 ;
        RECT 63.000 79.800 63.400 80.200 ;
        RECT 59.800 79.100 60.200 79.200 ;
        RECT 60.600 79.100 61.000 79.200 ;
        RECT 58.200 78.800 59.300 79.100 ;
        RECT 59.800 78.800 61.000 79.100 ;
        RECT 55.800 77.800 56.200 78.200 ;
        RECT 58.200 77.800 58.600 78.200 ;
        RECT 55.800 77.200 56.100 77.800 ;
        RECT 58.200 77.200 58.500 77.800 ;
        RECT 59.000 77.200 59.300 78.800 ;
        RECT 61.400 77.800 61.800 78.200 ;
        RECT 55.800 76.800 56.200 77.200 ;
        RECT 58.200 76.800 58.600 77.200 ;
        RECT 59.000 76.800 59.400 77.200 ;
        RECT 53.400 75.800 53.800 76.200 ;
        RECT 50.200 74.800 50.600 75.200 ;
        RECT 53.400 73.200 53.700 75.800 ;
        RECT 54.200 75.100 54.600 75.200 ;
        RECT 55.000 75.100 55.400 75.200 ;
        RECT 54.200 74.800 55.400 75.100 ;
        RECT 60.600 74.800 61.000 75.200 ;
        RECT 60.600 74.200 60.900 74.800 ;
        RECT 60.600 73.800 61.000 74.200 ;
        RECT 38.200 72.800 38.600 73.200 ;
        RECT 42.200 72.800 42.600 73.200 ;
        RECT 43.800 73.100 44.200 73.200 ;
        RECT 44.600 73.100 45.000 73.200 ;
        RECT 43.800 72.800 45.000 73.100 ;
        RECT 45.400 72.800 45.800 73.200 ;
        RECT 52.600 72.800 53.000 73.200 ;
        RECT 53.400 72.800 53.800 73.200 ;
        RECT 35.000 71.800 35.400 72.200 ;
        RECT 35.800 71.800 36.200 72.200 ;
        RECT 35.000 70.200 35.300 71.800 ;
        RECT 34.200 69.800 34.600 70.200 ;
        RECT 35.000 69.800 35.400 70.200 ;
        RECT 34.200 69.200 34.500 69.800 ;
        RECT 35.800 69.200 36.100 71.800 ;
        RECT 38.200 70.200 38.500 72.800 ;
        RECT 45.400 72.200 45.700 72.800 ;
        RECT 44.600 71.800 45.000 72.200 ;
        RECT 45.400 71.800 45.800 72.200 ;
        RECT 39.800 71.100 40.200 71.200 ;
        RECT 39.000 70.800 40.200 71.100 ;
        RECT 36.600 69.800 37.000 70.200 ;
        RECT 38.200 69.800 38.600 70.200 ;
        RECT 36.600 69.200 36.900 69.800 ;
        RECT 30.200 68.800 30.600 69.200 ;
        RECT 31.000 68.800 31.400 69.200 ;
        RECT 31.800 68.800 32.200 69.200 ;
        RECT 34.200 68.800 34.600 69.200 ;
        RECT 35.800 68.800 36.200 69.200 ;
        RECT 36.600 68.800 37.000 69.200 ;
        RECT 31.000 68.200 31.300 68.800 ;
        RECT 38.200 68.200 38.500 69.800 ;
        RECT 39.000 69.200 39.300 70.800 ;
        RECT 44.600 69.200 44.900 71.800 ;
        RECT 52.600 69.200 52.900 72.800 ;
        RECT 53.400 69.200 53.700 72.800 ;
        RECT 60.600 71.800 61.000 72.200 ;
        RECT 57.400 70.800 57.800 71.200 ;
        RECT 39.000 68.800 39.400 69.200 ;
        RECT 44.600 68.800 45.000 69.200 ;
        RECT 45.400 68.800 45.800 69.200 ;
        RECT 52.600 68.800 53.000 69.200 ;
        RECT 53.400 68.800 53.800 69.200 ;
        RECT 55.800 68.800 56.200 69.200 ;
        RECT 45.400 68.200 45.700 68.800 ;
        RECT 28.600 67.800 29.000 68.200 ;
        RECT 31.000 67.800 31.400 68.200 ;
        RECT 38.200 67.800 38.600 68.200 ;
        RECT 45.400 67.800 45.800 68.200 ;
        RECT 28.600 67.200 28.900 67.800 ;
        RECT 55.800 67.200 56.100 68.800 ;
        RECT 57.400 67.200 57.700 70.800 ;
        RECT 60.600 68.200 60.900 71.800 ;
        RECT 61.400 69.200 61.700 77.800 ;
        RECT 63.000 76.200 63.300 79.800 ;
        RECT 64.600 79.200 64.900 83.800 ;
        RECT 64.600 78.800 65.000 79.200 ;
        RECT 63.000 75.800 63.400 76.200 ;
        RECT 62.200 74.800 62.600 75.200 ;
        RECT 62.200 73.200 62.500 74.800 ;
        RECT 62.200 72.800 62.600 73.200 ;
        RECT 61.400 68.800 61.800 69.200 ;
        RECT 58.200 67.800 58.600 68.200 ;
        RECT 60.600 68.100 61.000 68.200 ;
        RECT 59.800 67.800 61.000 68.100 ;
        RECT 27.800 66.800 28.200 67.200 ;
        RECT 28.600 66.800 29.000 67.200 ;
        RECT 42.200 66.800 42.600 67.200 ;
        RECT 50.200 66.800 50.600 67.200 ;
        RECT 55.800 66.800 56.200 67.200 ;
        RECT 57.400 66.800 57.800 67.200 ;
        RECT 19.000 66.100 19.400 66.200 ;
        RECT 19.800 66.100 20.200 66.200 ;
        RECT 19.000 65.800 20.200 66.100 ;
        RECT 20.600 65.800 21.000 66.200 ;
        RECT 22.200 65.800 22.600 66.200 ;
        RECT 23.800 65.800 24.200 66.200 ;
        RECT 25.400 65.800 25.800 66.200 ;
        RECT 27.000 65.800 27.400 66.200 ;
        RECT 27.000 65.200 27.300 65.800 ;
        RECT 15.000 64.800 15.400 65.200 ;
        RECT 15.800 64.800 16.200 65.200 ;
        RECT 17.400 64.800 17.800 65.200 ;
        RECT 27.000 64.800 27.400 65.200 ;
        RECT 39.000 65.100 39.400 65.200 ;
        RECT 39.800 65.100 40.200 65.200 ;
        RECT 39.000 64.800 40.200 65.100 ;
        RECT 14.200 63.800 14.600 64.200 ;
        RECT 14.200 61.200 14.500 63.800 ;
        RECT 14.200 60.800 14.600 61.200 ;
        RECT 13.400 58.800 13.800 59.200 ;
        RECT 11.800 56.800 12.200 57.200 ;
        RECT 15.000 56.200 15.300 64.800 ;
        RECT 15.800 64.200 16.100 64.800 ;
        RECT 15.800 63.800 16.200 64.200 ;
        RECT 16.600 63.800 17.000 64.200 ;
        RECT 19.000 63.800 19.400 64.200 ;
        RECT 16.600 63.100 16.900 63.800 ;
        RECT 15.800 62.800 16.900 63.100 ;
        RECT 15.800 60.200 16.100 62.800 ;
        RECT 15.800 59.800 16.200 60.200 ;
        RECT 11.000 55.800 12.100 56.100 ;
        RECT 10.200 54.800 10.600 55.200 ;
        RECT 11.000 54.800 11.400 55.200 ;
        RECT 7.800 52.800 8.200 53.200 ;
        RECT 6.200 48.800 6.600 49.200 ;
        RECT 7.000 48.800 7.400 49.200 ;
        RECT 7.800 48.200 8.100 52.800 ;
        RECT 8.600 51.800 9.000 52.200 ;
        RECT 7.800 47.800 8.200 48.200 ;
        RECT 8.600 47.200 8.900 51.800 ;
        RECT 10.200 49.200 10.500 54.800 ;
        RECT 11.000 54.200 11.300 54.800 ;
        RECT 11.000 53.800 11.400 54.200 ;
        RECT 9.400 48.800 9.800 49.200 ;
        RECT 10.200 48.800 10.600 49.200 ;
        RECT 9.400 47.200 9.700 48.800 ;
        RECT 11.000 47.800 11.400 48.200 ;
        RECT 2.200 46.600 2.600 47.000 ;
        RECT 3.000 46.800 3.400 47.200 ;
        RECT 3.800 46.800 4.200 47.200 ;
        RECT 5.400 46.800 5.800 47.200 ;
        RECT 8.600 46.800 9.000 47.200 ;
        RECT 9.400 46.800 9.800 47.200 ;
        RECT 3.000 45.200 3.300 46.800 ;
        RECT 5.400 46.200 5.700 46.800 ;
        RECT 5.400 45.800 5.800 46.200 ;
        RECT 7.000 46.100 7.400 46.200 ;
        RECT 7.800 46.100 8.200 46.200 ;
        RECT 7.000 45.800 8.200 46.100 ;
        RECT 1.400 44.800 2.500 45.100 ;
        RECT 3.000 44.800 3.400 45.200 ;
        RECT 5.400 45.100 5.800 45.200 ;
        RECT 6.200 45.100 6.600 45.200 ;
        RECT 5.400 44.800 6.600 45.100 ;
        RECT 8.600 44.800 9.000 45.200 ;
        RECT 0.600 41.800 1.000 42.200 ;
        RECT 0.600 36.200 0.900 41.800 ;
        RECT 2.200 39.200 2.500 44.800 ;
        RECT 7.800 43.800 8.200 44.200 ;
        RECT 7.800 39.200 8.100 43.800 ;
        RECT 8.600 42.200 8.900 44.800 ;
        RECT 8.600 41.800 9.000 42.200 ;
        RECT 2.200 38.800 2.600 39.200 ;
        RECT 7.800 38.800 8.200 39.200 ;
        RECT 7.800 37.100 8.200 37.200 ;
        RECT 8.600 37.100 9.000 37.200 ;
        RECT 7.800 36.800 9.000 37.100 ;
        RECT 0.600 35.800 1.000 36.200 ;
        RECT 7.000 35.800 7.400 36.200 ;
        RECT 7.000 35.200 7.300 35.800 ;
        RECT 2.200 35.100 2.600 35.200 ;
        RECT 3.000 35.100 3.400 35.200 ;
        RECT 2.200 34.800 3.400 35.100 ;
        RECT 3.800 35.100 4.200 35.200 ;
        RECT 4.600 35.100 5.000 35.200 ;
        RECT 3.800 34.800 5.000 35.100 ;
        RECT 7.000 34.800 7.400 35.200 ;
        RECT 7.800 35.100 8.200 35.200 ;
        RECT 8.600 35.100 9.000 35.200 ;
        RECT 7.800 34.800 9.000 35.100 ;
        RECT 3.000 34.100 3.400 34.200 ;
        RECT 3.800 34.100 4.200 34.200 ;
        RECT 3.000 33.800 4.200 34.100 ;
        RECT 4.600 33.800 5.000 34.200 ;
        RECT 5.400 33.800 5.800 34.200 ;
        RECT 6.200 33.800 6.600 34.200 ;
        RECT 4.600 31.200 4.900 33.800 ;
        RECT 5.400 33.200 5.700 33.800 ;
        RECT 6.200 33.200 6.500 33.800 ;
        RECT 5.400 32.800 5.800 33.200 ;
        RECT 6.200 32.800 6.600 33.200 ;
        RECT 7.000 33.100 7.300 34.800 ;
        RECT 7.800 34.200 8.100 34.800 ;
        RECT 7.800 33.800 8.200 34.200 ;
        RECT 7.000 32.800 8.100 33.100 ;
        RECT 7.000 31.800 7.400 32.200 ;
        RECT 4.600 30.800 5.000 31.200 ;
        RECT 7.000 29.200 7.300 31.800 ;
        RECT 0.600 28.800 1.000 29.200 ;
        RECT 7.000 28.800 7.400 29.200 ;
        RECT 0.600 27.200 0.900 28.800 ;
        RECT 1.400 27.500 1.800 27.900 ;
        RECT 2.100 27.500 4.200 27.800 ;
        RECT 4.700 27.500 5.100 27.900 ;
        RECT 0.600 26.800 1.000 27.200 ;
        RECT 1.400 27.100 1.700 27.500 ;
        RECT 2.100 27.400 2.500 27.500 ;
        RECT 3.800 27.400 4.200 27.500 ;
        RECT 1.400 26.800 3.800 27.100 ;
        RECT 1.400 25.100 1.700 26.800 ;
        RECT 3.400 26.700 3.800 26.800 ;
        RECT 2.200 25.800 2.600 26.200 ;
        RECT 1.400 24.700 1.800 25.100 ;
        RECT 2.200 19.200 2.500 25.800 ;
        RECT 3.800 24.800 4.200 25.200 ;
        RECT 4.800 25.100 5.100 27.500 ;
        RECT 5.400 27.800 5.800 28.200 ;
        RECT 5.400 27.200 5.700 27.800 ;
        RECT 5.400 26.800 5.800 27.200 ;
        RECT 7.800 26.200 8.100 32.800 ;
        RECT 9.400 28.200 9.700 46.800 ;
        RECT 11.000 45.200 11.300 47.800 ;
        RECT 11.000 44.800 11.400 45.200 ;
        RECT 11.000 43.800 11.400 44.200 ;
        RECT 11.000 39.200 11.300 43.800 ;
        RECT 11.800 43.200 12.100 55.800 ;
        RECT 15.000 55.800 15.400 56.200 ;
        RECT 15.000 55.200 15.300 55.800 ;
        RECT 12.600 55.100 13.000 55.200 ;
        RECT 13.400 55.100 13.800 55.200 ;
        RECT 12.600 54.800 13.800 55.100 ;
        RECT 15.000 54.800 15.400 55.200 ;
        RECT 13.400 51.200 13.700 54.800 ;
        RECT 15.800 54.200 16.100 59.800 ;
        RECT 19.000 59.200 19.300 63.800 ;
        RECT 25.400 63.100 25.800 63.200 ;
        RECT 26.200 63.100 26.600 63.200 ;
        RECT 25.400 62.800 26.600 63.100 ;
        RECT 21.400 60.800 21.800 61.200 ;
        RECT 21.400 59.200 21.700 60.800 ;
        RECT 35.000 59.800 35.400 60.200 ;
        RECT 35.000 59.200 35.300 59.800 ;
        RECT 19.000 58.800 19.400 59.200 ;
        RECT 21.400 58.800 21.800 59.200 ;
        RECT 24.600 58.800 25.000 59.200 ;
        RECT 35.000 58.800 35.400 59.200 ;
        RECT 24.600 58.200 24.900 58.800 ;
        RECT 19.800 57.800 20.200 58.200 ;
        RECT 24.600 57.800 25.000 58.200 ;
        RECT 31.800 57.800 32.200 58.200 ;
        RECT 19.800 57.200 20.100 57.800 ;
        RECT 19.800 56.800 20.200 57.200 ;
        RECT 22.200 57.100 22.600 57.200 ;
        RECT 23.000 57.100 23.400 57.200 ;
        RECT 22.200 56.800 23.400 57.100 ;
        RECT 25.400 56.800 25.800 57.200 ;
        RECT 17.400 56.100 17.800 56.200 ;
        RECT 18.200 56.100 18.600 56.200 ;
        RECT 17.400 55.800 18.600 56.100 ;
        RECT 19.000 55.800 19.400 56.200 ;
        RECT 23.800 55.800 24.200 56.200 ;
        RECT 19.000 55.200 19.300 55.800 ;
        RECT 19.000 54.800 19.400 55.200 ;
        RECT 22.200 55.100 22.600 55.200 ;
        RECT 23.000 55.100 23.400 55.200 ;
        RECT 22.200 54.800 23.400 55.100 ;
        RECT 23.800 54.200 24.100 55.800 ;
        RECT 14.200 54.100 14.600 54.200 ;
        RECT 15.000 54.100 15.400 54.200 ;
        RECT 14.200 53.800 15.400 54.100 ;
        RECT 15.800 53.800 16.200 54.200 ;
        RECT 17.400 53.800 17.800 54.200 ;
        RECT 23.800 53.800 24.200 54.200 ;
        RECT 24.600 53.800 25.000 54.200 ;
        RECT 25.400 54.100 25.700 56.800 ;
        RECT 31.800 56.200 32.100 57.800 ;
        RECT 32.600 56.800 33.000 57.200 ;
        RECT 35.800 57.100 36.200 57.200 ;
        RECT 36.600 57.100 37.000 57.200 ;
        RECT 35.800 56.800 37.000 57.100 ;
        RECT 37.400 56.800 37.800 57.200 ;
        RECT 27.000 56.100 27.400 56.200 ;
        RECT 27.000 55.800 28.100 56.100 ;
        RECT 26.200 55.100 26.600 55.200 ;
        RECT 26.200 54.800 27.300 55.100 ;
        RECT 25.400 53.800 26.500 54.100 ;
        RECT 17.400 53.200 17.700 53.800 ;
        RECT 17.400 52.800 17.800 53.200 ;
        RECT 17.400 52.200 17.700 52.800 ;
        RECT 15.800 51.800 16.200 52.200 ;
        RECT 16.600 51.800 17.000 52.200 ;
        RECT 17.400 51.800 17.800 52.200 ;
        RECT 13.400 50.800 13.800 51.200 ;
        RECT 14.200 46.800 14.600 47.200 ;
        RECT 14.200 46.200 14.500 46.800 ;
        RECT 14.200 45.800 14.600 46.200 ;
        RECT 15.800 45.200 16.100 51.800 ;
        RECT 16.600 50.200 16.900 51.800 ;
        RECT 16.600 49.800 17.000 50.200 ;
        RECT 23.800 49.800 24.200 50.200 ;
        RECT 18.200 48.800 18.600 49.200 ;
        RECT 18.200 48.200 18.500 48.800 ;
        RECT 16.600 47.800 17.000 48.200 ;
        RECT 18.200 47.800 18.600 48.200 ;
        RECT 19.000 47.800 19.400 48.200 ;
        RECT 16.600 47.200 16.900 47.800 ;
        RECT 19.000 47.200 19.300 47.800 ;
        RECT 19.800 47.500 20.200 47.900 ;
        RECT 20.500 47.500 22.600 47.800 ;
        RECT 23.100 47.500 23.500 47.900 ;
        RECT 16.600 46.800 17.000 47.200 ;
        RECT 19.000 46.800 19.400 47.200 ;
        RECT 19.800 47.100 20.100 47.500 ;
        RECT 20.500 47.400 20.900 47.500 ;
        RECT 22.200 47.400 22.600 47.500 ;
        RECT 19.800 46.800 22.200 47.100 ;
        RECT 19.000 46.200 19.300 46.800 ;
        RECT 16.600 46.100 17.000 46.200 ;
        RECT 17.400 46.100 17.800 46.200 ;
        RECT 16.600 45.800 17.800 46.100 ;
        RECT 19.000 45.800 19.400 46.200 ;
        RECT 14.200 44.800 14.600 45.200 ;
        RECT 15.800 44.800 16.200 45.200 ;
        RECT 14.200 44.200 14.500 44.800 ;
        RECT 14.200 43.800 14.600 44.200 ;
        RECT 11.800 42.800 12.200 43.200 ;
        RECT 14.200 42.800 14.600 43.200 ;
        RECT 14.200 39.200 14.500 42.800 ;
        RECT 11.000 38.800 11.400 39.200 ;
        RECT 14.200 38.800 14.600 39.200 ;
        RECT 15.000 37.800 15.400 38.200 ;
        RECT 15.000 37.200 15.300 37.800 ;
        RECT 12.600 36.800 13.000 37.200 ;
        RECT 15.000 36.800 15.400 37.200 ;
        RECT 12.600 36.200 12.900 36.800 ;
        RECT 12.600 35.800 13.000 36.200 ;
        RECT 13.400 35.800 13.800 36.200 ;
        RECT 11.000 34.800 11.400 35.200 ;
        RECT 10.200 33.800 10.600 34.200 ;
        RECT 10.200 33.200 10.500 33.800 ;
        RECT 10.200 32.800 10.600 33.200 ;
        RECT 10.200 30.800 10.600 31.200 ;
        RECT 9.400 27.800 9.800 28.200 ;
        RECT 10.200 27.200 10.500 30.800 ;
        RECT 11.000 29.200 11.300 34.800 ;
        RECT 13.400 32.200 13.700 35.800 ;
        RECT 14.200 34.800 14.600 35.200 ;
        RECT 14.200 32.200 14.500 34.800 ;
        RECT 15.800 34.200 16.100 44.800 ;
        RECT 19.000 39.200 19.300 45.800 ;
        RECT 19.800 45.100 20.100 46.800 ;
        RECT 21.800 46.700 22.200 46.800 ;
        RECT 23.200 45.100 23.500 47.500 ;
        RECT 19.800 44.700 20.200 45.100 ;
        RECT 23.100 44.700 23.500 45.100 ;
        RECT 23.800 47.200 24.100 49.800 ;
        RECT 24.600 48.200 24.900 53.800 ;
        RECT 25.400 50.800 25.800 51.200 ;
        RECT 25.400 49.200 25.700 50.800 ;
        RECT 25.400 48.800 25.800 49.200 ;
        RECT 24.600 47.800 25.000 48.200 ;
        RECT 26.200 47.200 26.500 53.800 ;
        RECT 27.000 48.200 27.300 54.800 ;
        RECT 27.800 53.200 28.100 55.800 ;
        RECT 31.000 55.800 31.400 56.200 ;
        RECT 31.800 55.800 32.200 56.200 ;
        RECT 29.400 55.100 29.800 55.200 ;
        RECT 30.200 55.100 30.600 55.200 ;
        RECT 29.400 54.800 30.600 55.100 ;
        RECT 31.000 54.200 31.300 55.800 ;
        RECT 31.800 54.800 32.200 55.200 ;
        RECT 29.400 53.800 29.800 54.200 ;
        RECT 31.000 53.800 31.400 54.200 ;
        RECT 27.800 53.100 28.200 53.200 ;
        RECT 28.600 53.100 29.000 53.200 ;
        RECT 27.800 52.800 29.000 53.100 ;
        RECT 29.400 52.200 29.700 53.800 ;
        RECT 27.800 52.100 28.200 52.200 ;
        RECT 28.600 52.100 29.000 52.200 ;
        RECT 27.800 51.800 29.000 52.100 ;
        RECT 29.400 51.800 29.800 52.200 ;
        RECT 27.000 47.800 27.400 48.200 ;
        RECT 23.800 46.800 24.200 47.200 ;
        RECT 26.200 46.800 26.600 47.200 ;
        RECT 20.600 41.800 21.000 42.200 ;
        RECT 21.400 41.800 21.800 42.200 ;
        RECT 20.600 39.200 20.900 41.800 ;
        RECT 19.000 38.800 19.400 39.200 ;
        RECT 20.600 38.800 21.000 39.200 ;
        RECT 21.400 38.200 21.700 41.800 ;
        RECT 21.400 37.800 21.800 38.200 ;
        RECT 18.200 36.800 18.600 37.200 ;
        RECT 20.600 37.100 21.000 37.200 ;
        RECT 21.400 37.100 21.800 37.200 ;
        RECT 23.800 37.100 24.100 46.800 ;
        RECT 27.000 46.200 27.300 47.800 ;
        RECT 31.800 47.200 32.100 54.800 ;
        RECT 32.600 52.200 32.900 56.800 ;
        RECT 34.200 55.800 34.600 56.200 ;
        RECT 34.200 53.200 34.500 55.800 ;
        RECT 35.000 55.100 35.400 55.200 ;
        RECT 35.800 55.100 36.200 55.200 ;
        RECT 35.000 54.800 36.200 55.100 ;
        RECT 37.400 54.200 37.700 56.800 ;
        RECT 39.800 55.200 40.100 64.800 ;
        RECT 42.200 63.200 42.500 66.800 ;
        RECT 43.000 65.800 43.400 66.200 ;
        RECT 42.200 62.800 42.600 63.200 ;
        RECT 42.200 55.200 42.500 62.800 ;
        RECT 43.000 55.200 43.300 65.800 ;
        RECT 45.400 64.800 45.800 65.200 ;
        RECT 44.600 61.800 45.000 62.200 ;
        RECT 44.600 55.200 44.900 61.800 ;
        RECT 45.400 59.200 45.700 64.800 ;
        RECT 50.200 59.200 50.500 66.800 ;
        RECT 58.200 66.200 58.500 67.800 ;
        RECT 59.800 67.200 60.100 67.800 ;
        RECT 59.800 66.800 60.200 67.200 ;
        RECT 60.600 66.800 61.000 67.200 ;
        RECT 51.000 65.800 51.400 66.200 ;
        RECT 56.600 65.800 57.000 66.200 ;
        RECT 58.200 65.800 58.600 66.200 ;
        RECT 45.400 58.800 45.800 59.200 ;
        RECT 48.600 59.100 49.000 59.200 ;
        RECT 49.400 59.100 49.800 59.200 ;
        RECT 48.600 58.800 49.800 59.100 ;
        RECT 50.200 58.800 50.600 59.200 ;
        RECT 51.000 55.200 51.300 65.800 ;
        RECT 52.600 64.800 53.000 65.200 ;
        RECT 38.200 54.800 38.600 55.200 ;
        RECT 39.000 54.800 39.400 55.200 ;
        RECT 39.800 54.800 40.200 55.200 ;
        RECT 40.600 55.100 41.000 55.200 ;
        RECT 41.400 55.100 41.800 55.200 ;
        RECT 40.600 54.800 41.800 55.100 ;
        RECT 42.200 54.800 42.600 55.200 ;
        RECT 43.000 54.800 43.400 55.200 ;
        RECT 44.600 54.800 45.000 55.200 ;
        RECT 45.400 54.800 45.800 55.200 ;
        RECT 51.000 54.800 51.400 55.200 ;
        RECT 37.400 53.800 37.800 54.200 ;
        RECT 34.200 52.800 34.600 53.200 ;
        RECT 32.600 51.800 33.000 52.200 ;
        RECT 37.400 51.800 37.800 52.200 ;
        RECT 37.400 49.200 37.700 51.800 ;
        RECT 37.400 48.800 37.800 49.200 ;
        RECT 38.200 48.200 38.500 54.800 ;
        RECT 39.000 54.200 39.300 54.800 ;
        RECT 39.000 53.800 39.400 54.200 ;
        RECT 41.400 53.800 41.800 54.200 ;
        RECT 41.400 53.100 41.700 53.800 ;
        RECT 42.200 53.100 42.600 53.200 ;
        RECT 41.400 52.800 42.600 53.100 ;
        RECT 44.600 52.100 44.900 54.800 ;
        RECT 45.400 53.200 45.700 54.800 ;
        RECT 47.000 53.800 47.400 54.200 ;
        RECT 51.000 53.800 51.400 54.200 ;
        RECT 45.400 52.800 45.800 53.200 ;
        RECT 46.200 52.800 46.600 53.200 ;
        RECT 46.200 52.200 46.500 52.800 ;
        RECT 44.600 51.800 45.700 52.100 ;
        RECT 46.200 51.800 46.600 52.200 ;
        RECT 35.800 47.800 36.200 48.200 ;
        RECT 38.200 47.800 38.600 48.200 ;
        RECT 40.600 47.800 41.000 48.200 ;
        RECT 42.200 47.800 42.600 48.200 ;
        RECT 43.000 48.100 43.400 48.200 ;
        RECT 43.800 48.100 44.200 48.200 ;
        RECT 43.000 47.800 44.200 48.100 ;
        RECT 35.800 47.200 36.100 47.800 ;
        RECT 30.200 47.100 30.600 47.200 ;
        RECT 31.000 47.100 31.400 47.200 ;
        RECT 30.200 46.800 31.400 47.100 ;
        RECT 31.800 46.800 32.200 47.200 ;
        RECT 34.200 46.800 34.600 47.200 ;
        RECT 35.800 46.800 36.200 47.200 ;
        RECT 39.800 46.800 40.200 47.200 ;
        RECT 27.000 45.800 27.400 46.200 ;
        RECT 29.400 46.100 29.800 46.200 ;
        RECT 30.200 46.100 30.600 46.200 ;
        RECT 29.400 45.800 30.600 46.100 ;
        RECT 34.200 45.200 34.500 46.800 ;
        RECT 39.800 46.200 40.100 46.800 ;
        RECT 40.600 46.200 40.900 47.800 ;
        RECT 35.000 45.800 35.400 46.200 ;
        RECT 38.200 46.100 38.600 46.200 ;
        RECT 39.000 46.100 39.400 46.200 ;
        RECT 38.200 45.800 39.400 46.100 ;
        RECT 39.800 45.800 40.200 46.200 ;
        RECT 40.600 45.800 41.000 46.200 ;
        RECT 27.800 44.800 28.200 45.200 ;
        RECT 31.000 44.800 31.400 45.200 ;
        RECT 34.200 44.800 34.600 45.200 ;
        RECT 27.800 44.200 28.100 44.800 ;
        RECT 31.000 44.200 31.300 44.800 ;
        RECT 27.800 43.800 28.200 44.200 ;
        RECT 31.000 43.800 31.400 44.200 ;
        RECT 31.000 39.200 31.300 43.800 ;
        RECT 34.200 42.800 34.600 43.200 ;
        RECT 34.200 39.200 34.500 42.800 ;
        RECT 20.600 36.800 21.800 37.100 ;
        RECT 23.000 36.800 24.100 37.100 ;
        RECT 27.800 38.800 28.200 39.200 ;
        RECT 31.000 38.800 31.400 39.200 ;
        RECT 34.200 38.800 34.600 39.200 ;
        RECT 16.600 34.800 17.000 35.200 ;
        RECT 16.600 34.200 16.900 34.800 ;
        RECT 18.200 34.200 18.500 36.800 ;
        RECT 19.800 35.800 20.200 36.200 ;
        RECT 15.000 33.800 15.400 34.200 ;
        RECT 15.800 33.800 16.200 34.200 ;
        RECT 16.600 33.800 17.000 34.200 ;
        RECT 18.200 33.800 18.600 34.200 ;
        RECT 13.400 31.800 13.800 32.200 ;
        RECT 14.200 31.800 14.600 32.200 ;
        RECT 15.000 29.200 15.300 33.800 ;
        RECT 15.800 29.200 16.100 33.800 ;
        RECT 16.600 33.100 17.000 33.200 ;
        RECT 17.400 33.100 17.800 33.200 ;
        RECT 16.600 32.800 17.800 33.100 ;
        RECT 11.000 28.800 11.400 29.200 ;
        RECT 15.000 28.800 15.400 29.200 ;
        RECT 15.800 28.800 16.200 29.200 ;
        RECT 11.800 27.800 12.200 28.200 ;
        RECT 18.200 28.100 18.500 33.800 ;
        RECT 19.000 31.800 19.400 32.200 ;
        RECT 19.000 29.200 19.300 31.800 ;
        RECT 19.000 28.800 19.400 29.200 ;
        RECT 18.200 27.800 19.300 28.100 ;
        RECT 10.200 26.800 10.600 27.200 ;
        RECT 7.000 26.100 7.400 26.200 ;
        RECT 7.800 26.100 8.200 26.200 ;
        RECT 7.000 25.800 8.200 26.100 ;
        RECT 8.600 26.100 9.000 26.200 ;
        RECT 9.400 26.100 9.800 26.200 ;
        RECT 8.600 25.800 9.800 26.100 ;
        RECT 3.800 24.200 4.100 24.800 ;
        RECT 4.700 24.700 5.100 25.100 ;
        RECT 7.800 25.100 8.200 25.200 ;
        RECT 8.600 25.100 9.000 25.200 ;
        RECT 7.800 24.800 9.000 25.100 ;
        RECT 10.200 24.200 10.500 26.800 ;
        RECT 11.800 25.200 12.100 27.800 ;
        RECT 13.400 27.100 13.800 27.200 ;
        RECT 14.200 27.100 14.600 27.200 ;
        RECT 13.400 26.800 14.600 27.100 ;
        RECT 15.800 26.800 16.200 27.200 ;
        RECT 17.400 26.800 17.800 27.200 ;
        RECT 11.800 24.800 12.200 25.200 ;
        RECT 15.800 24.200 16.100 26.800 ;
        RECT 16.600 25.800 17.000 26.200 ;
        RECT 16.600 25.200 16.900 25.800 ;
        RECT 17.400 25.200 17.700 26.800 ;
        RECT 18.200 25.800 18.600 26.200 ;
        RECT 16.600 24.800 17.000 25.200 ;
        RECT 17.400 24.800 17.800 25.200 ;
        RECT 3.800 23.800 4.200 24.200 ;
        RECT 8.600 23.800 9.000 24.200 ;
        RECT 10.200 23.800 10.600 24.200 ;
        RECT 15.800 23.800 16.200 24.200 ;
        RECT 8.600 19.200 8.900 23.800 ;
        RECT 18.200 19.200 18.500 25.800 ;
        RECT 19.000 24.200 19.300 27.800 ;
        RECT 19.800 26.200 20.100 35.800 ;
        RECT 23.000 35.200 23.300 36.800 ;
        RECT 23.900 35.900 24.300 36.300 ;
        RECT 24.600 36.100 25.000 36.200 ;
        RECT 25.400 36.100 25.800 36.200 ;
        RECT 20.600 35.100 21.000 35.200 ;
        RECT 21.400 35.100 21.800 35.200 ;
        RECT 20.600 34.800 21.800 35.100 ;
        RECT 23.000 34.800 23.400 35.200 ;
        RECT 20.600 33.200 20.900 34.800 ;
        RECT 23.000 34.200 23.300 34.800 ;
        RECT 23.000 33.800 23.400 34.200 ;
        RECT 23.900 33.500 24.200 35.900 ;
        RECT 24.600 35.800 25.800 36.100 ;
        RECT 27.000 35.900 27.400 36.300 ;
        RECT 24.500 34.900 24.900 35.300 ;
        RECT 24.600 34.200 24.900 34.900 ;
        RECT 27.100 34.200 27.400 35.900 ;
        RECT 24.600 33.900 27.400 34.200 ;
        RECT 24.600 33.500 25.000 33.600 ;
        RECT 26.300 33.500 26.700 33.600 ;
        RECT 27.100 33.500 27.400 33.900 ;
        RECT 27.800 34.200 28.100 38.800 ;
        RECT 35.000 37.200 35.300 45.800 ;
        RECT 36.600 44.800 37.000 45.200 ;
        RECT 40.600 44.800 41.000 45.200 ;
        RECT 36.600 39.200 36.900 44.800 ;
        RECT 40.600 44.200 40.900 44.800 ;
        RECT 42.200 44.200 42.500 47.800 ;
        RECT 43.000 47.100 43.400 47.200 ;
        RECT 43.800 47.100 44.200 47.200 ;
        RECT 43.000 46.800 44.200 47.100 ;
        RECT 45.400 46.200 45.700 51.800 ;
        RECT 47.000 50.200 47.300 53.800 ;
        RECT 51.000 53.200 51.300 53.800 ;
        RECT 52.600 53.200 52.900 64.800 ;
        RECT 55.800 62.800 56.200 63.200 ;
        RECT 55.800 59.200 56.100 62.800 ;
        RECT 55.800 58.800 56.200 59.200 ;
        RECT 56.600 55.200 56.900 65.800 ;
        RECT 60.600 61.200 60.900 66.800 ;
        RECT 60.600 60.800 61.000 61.200 ;
        RECT 61.400 59.200 61.700 68.800 ;
        RECT 63.000 68.200 63.300 75.800 ;
        RECT 64.600 74.800 65.000 75.200 ;
        RECT 64.600 69.200 64.900 74.800 ;
        RECT 65.400 71.200 65.700 85.800 ;
        RECT 66.200 85.200 66.500 86.800 ;
        RECT 66.200 84.800 66.600 85.200 ;
        RECT 67.000 85.100 67.400 85.200 ;
        RECT 67.000 84.800 68.100 85.100 ;
        RECT 66.200 75.200 66.500 84.800 ;
        RECT 67.000 83.800 67.400 84.200 ;
        RECT 67.000 79.200 67.300 83.800 ;
        RECT 67.000 78.800 67.400 79.200 ;
        RECT 67.800 77.100 68.100 84.800 ;
        RECT 68.600 84.200 68.900 93.800 ;
        RECT 69.400 95.200 69.700 95.800 ;
        RECT 74.200 95.200 74.500 95.800 ;
        RECT 77.400 95.200 77.700 97.800 ;
        RECT 87.000 97.200 87.300 101.800 ;
        RECT 78.200 97.100 78.600 97.200 ;
        RECT 79.000 97.100 79.400 97.200 ;
        RECT 78.200 96.800 79.400 97.100 ;
        RECT 87.000 96.800 87.400 97.200 ;
        RECT 81.400 95.800 81.800 96.200 ;
        RECT 87.000 95.800 87.400 96.200 ;
        RECT 81.400 95.200 81.700 95.800 ;
        RECT 87.000 95.200 87.300 95.800 ;
        RECT 69.400 94.800 69.800 95.200 ;
        RECT 71.800 94.800 72.200 95.200 ;
        RECT 74.200 94.800 74.600 95.200 ;
        RECT 75.000 95.100 75.400 95.200 ;
        RECT 75.800 95.100 76.200 95.200 ;
        RECT 75.000 94.800 76.200 95.100 ;
        RECT 76.600 94.800 77.000 95.200 ;
        RECT 77.400 94.800 77.800 95.200 ;
        RECT 79.000 94.800 79.400 95.200 ;
        RECT 79.800 95.100 80.200 95.200 ;
        RECT 80.600 95.100 81.000 95.200 ;
        RECT 79.800 94.800 81.000 95.100 ;
        RECT 81.400 94.800 81.800 95.200 ;
        RECT 83.000 94.800 83.400 95.200 ;
        RECT 87.000 94.800 87.400 95.200 ;
        RECT 69.400 91.200 69.700 94.800 ;
        RECT 71.800 94.200 72.100 94.800 ;
        RECT 71.800 93.800 72.200 94.200 ;
        RECT 72.600 94.100 73.000 94.200 ;
        RECT 73.400 94.100 73.800 94.200 ;
        RECT 72.600 93.800 73.800 94.100 ;
        RECT 75.000 93.800 75.400 94.200 ;
        RECT 75.000 93.200 75.300 93.800 ;
        RECT 71.800 93.100 72.200 93.200 ;
        RECT 72.600 93.100 73.000 93.200 ;
        RECT 71.800 92.800 73.000 93.100 ;
        RECT 75.000 92.800 75.400 93.200 ;
        RECT 76.600 92.200 76.900 94.800 ;
        RECT 77.400 94.100 77.800 94.200 ;
        RECT 78.200 94.100 78.600 94.200 ;
        RECT 77.400 93.800 78.600 94.100 ;
        RECT 71.000 91.800 71.400 92.200 ;
        RECT 76.600 91.800 77.000 92.200 ;
        RECT 69.400 90.800 69.800 91.200 ;
        RECT 70.200 86.800 70.600 87.200 ;
        RECT 69.400 85.800 69.800 86.200 ;
        RECT 68.600 83.800 69.000 84.200 ;
        RECT 68.600 77.100 69.000 77.200 ;
        RECT 67.800 76.800 69.000 77.100 ;
        RECT 68.600 76.200 68.900 76.800 ;
        RECT 68.600 75.800 69.000 76.200 ;
        RECT 66.200 74.800 66.600 75.200 ;
        RECT 69.400 75.100 69.700 85.800 ;
        RECT 70.200 79.200 70.500 86.800 ;
        RECT 70.200 78.800 70.600 79.200 ;
        RECT 68.600 74.800 69.700 75.100 ;
        RECT 71.000 75.200 71.300 91.800 ;
        RECT 71.800 90.800 72.200 91.200 ;
        RECT 71.800 87.200 72.100 90.800 ;
        RECT 79.000 89.200 79.300 94.800 ;
        RECT 80.600 93.800 81.000 94.200 ;
        RECT 80.600 92.200 80.900 93.800 ;
        RECT 80.600 91.800 81.000 92.200 ;
        RECT 81.400 90.200 81.700 94.800 ;
        RECT 83.000 93.200 83.300 94.800 ;
        RECT 83.800 93.800 84.200 94.200 ;
        RECT 83.000 92.800 83.400 93.200 ;
        RECT 83.800 92.200 84.100 93.800 ;
        RECT 83.800 91.800 84.200 92.200 ;
        RECT 84.600 91.800 85.000 92.200 ;
        RECT 81.400 89.800 81.800 90.200 ;
        RECT 83.800 89.200 84.100 91.800 ;
        RECT 84.600 89.200 84.900 91.800 ;
        RECT 87.800 89.200 88.100 101.800 ;
        RECT 91.000 99.200 91.300 103.800 ;
        RECT 99.000 101.200 99.300 107.800 ;
        RECT 102.200 105.800 102.600 106.200 ;
        RECT 99.000 100.800 99.400 101.200 ;
        RECT 91.000 98.800 91.400 99.200 ;
        RECT 97.400 98.800 97.800 99.200 ;
        RECT 89.400 97.800 89.800 98.200 ;
        RECT 96.600 97.800 97.000 98.200 ;
        RECT 89.400 96.200 89.700 97.800 ;
        RECT 96.600 97.200 96.900 97.800 ;
        RECT 95.000 97.100 95.400 97.200 ;
        RECT 95.800 97.100 96.200 97.200 ;
        RECT 95.000 96.800 96.200 97.100 ;
        RECT 96.600 96.800 97.000 97.200 ;
        RECT 97.400 96.200 97.700 98.800 ;
        RECT 99.000 96.800 99.400 97.200 ;
        RECT 99.000 96.200 99.300 96.800 ;
        RECT 102.200 96.200 102.500 105.800 ;
        RECT 107.000 102.100 107.400 108.900 ;
        RECT 107.800 102.100 108.200 108.900 ;
        RECT 108.600 103.100 109.000 108.900 ;
        RECT 109.400 106.800 109.800 107.200 ;
        RECT 106.200 100.800 106.600 101.200 ;
        RECT 106.200 99.200 106.500 100.800 ;
        RECT 109.400 99.200 109.700 106.800 ;
        RECT 110.200 103.100 110.600 108.900 ;
        RECT 111.800 103.100 112.200 108.900 ;
        RECT 112.600 102.100 113.000 108.900 ;
        RECT 113.400 102.100 113.800 108.900 ;
        RECT 114.200 102.100 114.600 108.900 ;
        RECT 120.600 108.100 121.000 108.200 ;
        RECT 121.400 108.100 121.800 108.200 ;
        RECT 120.600 107.800 121.800 108.100 ;
        RECT 115.000 105.800 115.400 106.200 ;
        RECT 115.000 104.200 115.300 105.800 ;
        RECT 115.800 104.800 116.200 105.200 ;
        RECT 119.800 105.100 120.200 105.200 ;
        RECT 120.600 105.100 121.000 105.200 ;
        RECT 119.800 104.800 121.000 105.100 ;
        RECT 115.000 103.800 115.400 104.200 ;
        RECT 115.800 99.200 116.100 104.800 ;
        RECT 119.000 102.100 119.400 102.200 ;
        RECT 119.800 102.100 120.200 102.200 ;
        RECT 119.000 101.800 120.200 102.100 ;
        RECT 121.400 101.800 121.800 102.200 ;
        RECT 106.200 98.800 106.600 99.200 ;
        RECT 109.400 98.800 109.800 99.200 ;
        RECT 115.800 98.800 116.200 99.200 ;
        RECT 119.800 99.100 120.200 99.200 ;
        RECT 120.600 99.100 121.000 99.200 ;
        RECT 119.800 98.800 121.000 99.100 ;
        RECT 105.400 97.800 105.800 98.200 ;
        RECT 105.400 96.200 105.700 97.800 ;
        RECT 89.400 95.800 89.800 96.200 ;
        RECT 96.600 95.800 97.000 96.200 ;
        RECT 97.400 95.800 97.800 96.200 ;
        RECT 99.000 95.800 99.400 96.200 ;
        RECT 102.200 95.800 102.600 96.200 ;
        RECT 105.400 95.800 105.800 96.200 ;
        RECT 96.600 95.200 96.900 95.800 ;
        RECT 91.000 94.800 91.400 95.200 ;
        RECT 91.800 95.100 92.200 95.200 ;
        RECT 92.600 95.100 93.000 95.200 ;
        RECT 91.800 94.800 93.000 95.100 ;
        RECT 96.600 94.800 97.000 95.200 ;
        RECT 88.600 93.800 89.000 94.200 ;
        RECT 88.600 90.200 88.900 93.800 ;
        RECT 91.000 92.200 91.300 94.800 ;
        RECT 91.800 94.100 92.200 94.200 ;
        RECT 92.600 94.100 93.000 94.200 ;
        RECT 91.800 93.800 93.000 94.100 ;
        RECT 96.600 93.800 97.000 94.200 ;
        RECT 92.600 92.800 93.000 93.200 ;
        RECT 93.400 93.100 93.800 93.200 ;
        RECT 94.200 93.100 94.600 93.200 ;
        RECT 93.400 92.800 94.600 93.100 ;
        RECT 91.000 91.800 91.400 92.200 ;
        RECT 88.600 89.800 89.000 90.200 ;
        RECT 92.600 90.100 92.900 92.800 ;
        RECT 91.800 89.800 92.900 90.100 ;
        RECT 73.400 89.100 73.800 89.200 ;
        RECT 74.200 89.100 74.600 89.200 ;
        RECT 73.400 88.800 74.600 89.100 ;
        RECT 79.000 88.800 79.400 89.200 ;
        RECT 83.800 88.800 84.200 89.200 ;
        RECT 84.600 88.800 85.000 89.200 ;
        RECT 87.000 88.800 87.400 89.200 ;
        RECT 87.800 88.800 88.200 89.200 ;
        RECT 87.000 88.200 87.300 88.800 ;
        RECT 91.800 88.200 92.100 89.800 ;
        RECT 92.600 89.100 93.000 89.200 ;
        RECT 93.400 89.100 93.800 89.200 ;
        RECT 92.600 88.800 93.800 89.100 ;
        RECT 76.600 87.500 77.000 87.900 ;
        RECT 79.700 87.800 80.100 87.900 ;
        RECT 77.300 87.500 80.100 87.800 ;
        RECT 71.800 86.800 72.200 87.200 ;
        RECT 75.800 86.800 76.200 87.200 ;
        RECT 76.600 87.100 76.900 87.500 ;
        RECT 77.300 87.400 77.700 87.500 ;
        RECT 79.000 87.400 79.400 87.500 ;
        RECT 76.600 86.800 79.400 87.100 ;
        RECT 75.800 86.200 76.100 86.800 ;
        RECT 75.800 85.800 76.200 86.200 ;
        RECT 72.600 84.800 73.000 85.200 ;
        RECT 72.600 80.200 72.900 84.800 ;
        RECT 75.800 81.200 76.100 85.800 ;
        RECT 76.600 85.100 76.900 86.800 ;
        RECT 79.100 86.100 79.400 86.800 ;
        RECT 79.100 85.700 79.500 86.100 ;
        RECT 79.800 85.100 80.100 87.500 ;
        RECT 87.000 87.800 87.400 88.200 ;
        RECT 91.800 87.800 92.200 88.200 ;
        RECT 94.200 88.100 94.600 88.200 ;
        RECT 95.000 88.100 95.400 88.200 ;
        RECT 94.200 87.800 95.400 88.100 ;
        RECT 76.600 84.700 77.000 85.100 ;
        RECT 79.700 84.700 80.100 85.100 ;
        RECT 80.600 86.800 81.000 87.200 ;
        RECT 73.400 80.800 73.800 81.200 ;
        RECT 75.800 80.800 76.200 81.200 ;
        RECT 72.600 79.800 73.000 80.200 ;
        RECT 71.800 79.100 72.200 79.200 ;
        RECT 72.600 79.100 73.000 79.200 ;
        RECT 71.800 78.800 73.000 79.100 ;
        RECT 71.000 74.800 71.400 75.200 ;
        RECT 72.600 74.800 73.000 75.200 ;
        RECT 66.200 73.800 66.600 74.200 ;
        RECT 65.400 70.800 65.800 71.200 ;
        RECT 66.200 69.200 66.500 73.800 ;
        RECT 68.600 72.200 68.900 74.800 ;
        RECT 69.400 72.800 69.800 73.200 ;
        RECT 69.400 72.200 69.700 72.800 ;
        RECT 68.600 71.800 69.000 72.200 ;
        RECT 69.400 71.800 69.800 72.200 ;
        RECT 71.000 69.200 71.300 74.800 ;
        RECT 72.600 74.200 72.900 74.800 ;
        RECT 71.800 73.800 72.200 74.200 ;
        RECT 72.600 73.800 73.000 74.200 ;
        RECT 71.800 72.200 72.100 73.800 ;
        RECT 71.800 71.800 72.200 72.200 ;
        RECT 64.600 68.800 65.000 69.200 ;
        RECT 66.200 68.800 66.600 69.200 ;
        RECT 67.800 69.100 68.200 69.200 ;
        RECT 68.600 69.100 69.000 69.200 ;
        RECT 67.800 68.800 69.000 69.100 ;
        RECT 71.000 68.800 71.400 69.200 ;
        RECT 71.000 68.200 71.300 68.800 ;
        RECT 63.000 67.800 63.400 68.200 ;
        RECT 63.800 68.100 64.200 68.200 ;
        RECT 64.600 68.100 65.000 68.200 ;
        RECT 63.800 67.800 65.000 68.100 ;
        RECT 69.400 68.100 69.800 68.200 ;
        RECT 70.200 68.100 70.600 68.200 ;
        RECT 69.400 67.800 70.600 68.100 ;
        RECT 71.000 67.800 71.400 68.200 ;
        RECT 65.400 66.800 65.800 67.200 ;
        RECT 63.000 66.100 63.400 66.200 ;
        RECT 63.800 66.100 64.200 66.200 ;
        RECT 63.000 65.800 64.200 66.100 ;
        RECT 63.800 62.800 64.200 63.200 ;
        RECT 63.800 59.200 64.100 62.800 ;
        RECT 57.400 59.100 57.800 59.200 ;
        RECT 58.200 59.100 58.600 59.200 ;
        RECT 57.400 58.800 58.600 59.100 ;
        RECT 61.400 58.800 61.800 59.200 ;
        RECT 63.800 58.800 64.200 59.200 ;
        RECT 63.000 57.800 63.400 58.200 ;
        RECT 53.400 55.100 53.800 55.200 ;
        RECT 54.200 55.100 54.600 55.200 ;
        RECT 53.400 54.800 54.600 55.100 ;
        RECT 56.600 54.800 57.000 55.200 ;
        RECT 59.800 55.100 60.200 55.200 ;
        RECT 60.600 55.100 61.000 55.200 ;
        RECT 59.800 54.800 61.000 55.100 ;
        RECT 51.000 52.800 51.400 53.200 ;
        RECT 51.800 52.800 52.200 53.200 ;
        RECT 52.600 52.800 53.000 53.200 ;
        RECT 53.400 52.800 53.800 53.200 ;
        RECT 55.000 52.800 55.400 53.200 ;
        RECT 56.600 53.100 56.900 54.800 ;
        RECT 63.000 54.200 63.300 57.800 ;
        RECT 64.600 54.800 65.000 55.200 ;
        RECT 60.600 53.800 61.000 54.200 ;
        RECT 63.000 53.800 63.400 54.200 ;
        RECT 60.600 53.200 60.900 53.800 ;
        RECT 57.400 53.100 57.800 53.200 ;
        RECT 56.600 52.800 57.800 53.100 ;
        RECT 60.600 52.800 61.000 53.200 ;
        RECT 51.800 52.200 52.100 52.800 ;
        RECT 51.800 51.800 52.200 52.200 ;
        RECT 47.000 49.800 47.400 50.200 ;
        RECT 53.400 49.200 53.700 52.800 ;
        RECT 55.000 52.200 55.300 52.800 ;
        RECT 55.000 51.800 55.400 52.200 ;
        RECT 55.000 50.200 55.300 51.800 ;
        RECT 54.200 49.800 54.600 50.200 ;
        RECT 55.000 49.800 55.400 50.200 ;
        RECT 53.400 48.800 53.800 49.200 ;
        RECT 46.200 47.800 46.600 48.200 ;
        RECT 49.400 48.100 49.800 48.200 ;
        RECT 50.200 48.100 50.600 48.200 ;
        RECT 49.400 47.800 50.600 48.100 ;
        RECT 51.000 47.800 51.400 48.200 ;
        RECT 46.200 47.200 46.500 47.800 ;
        RECT 46.200 46.800 46.600 47.200 ;
        RECT 47.800 46.800 48.200 47.200 ;
        RECT 48.600 47.100 49.000 47.200 ;
        RECT 49.400 47.100 49.800 47.200 ;
        RECT 48.600 46.800 49.800 47.100 ;
        RECT 47.800 46.200 48.100 46.800 ;
        RECT 51.000 46.200 51.300 47.800 ;
        RECT 54.200 47.200 54.500 49.800 ;
        RECT 57.400 49.200 57.700 52.800 ;
        RECT 63.800 51.800 64.200 52.200 ;
        RECT 61.400 49.800 61.800 50.200 ;
        RECT 63.000 49.800 63.400 50.200 ;
        RECT 61.400 49.200 61.700 49.800 ;
        RECT 57.400 48.800 57.800 49.200 ;
        RECT 61.400 48.800 61.800 49.200 ;
        RECT 54.200 46.800 54.600 47.200 ;
        RECT 55.000 46.800 55.400 47.200 ;
        RECT 55.800 46.800 56.200 47.200 ;
        RECT 57.400 47.100 57.800 47.200 ;
        RECT 58.200 47.100 58.600 47.200 ;
        RECT 57.400 46.800 58.600 47.100 ;
        RECT 59.000 46.800 59.400 47.200 ;
        RECT 60.600 47.100 61.000 47.200 ;
        RECT 61.400 47.100 61.800 47.200 ;
        RECT 60.600 46.800 61.800 47.100 ;
        RECT 45.400 46.100 45.800 46.200 ;
        RECT 46.200 46.100 46.600 46.200 ;
        RECT 45.400 45.800 46.600 46.100 ;
        RECT 47.800 45.800 48.200 46.200 ;
        RECT 51.000 45.800 51.400 46.200 ;
        RECT 52.600 45.800 53.000 46.200 ;
        RECT 40.600 43.800 41.000 44.200 ;
        RECT 42.200 43.800 42.600 44.200 ;
        RECT 36.600 38.800 37.000 39.200 ;
        RECT 39.800 38.800 40.200 39.200 ;
        RECT 39.800 38.200 40.100 38.800 ;
        RECT 39.800 37.800 40.200 38.200 ;
        RECT 35.000 36.800 35.400 37.200 ;
        RECT 41.400 37.100 41.800 37.200 ;
        RECT 42.200 37.100 42.600 37.200 ;
        RECT 41.400 36.800 42.600 37.100 ;
        RECT 27.800 33.800 28.200 34.200 ;
        RECT 23.900 33.200 26.700 33.500 ;
        RECT 20.600 32.800 21.000 33.200 ;
        RECT 23.900 33.100 24.300 33.200 ;
        RECT 27.000 33.100 27.400 33.500 ;
        RECT 31.800 33.100 32.200 33.200 ;
        RECT 32.600 33.100 33.000 33.200 ;
        RECT 31.800 32.800 33.000 33.100 ;
        RECT 28.600 31.800 29.000 32.200 ;
        RECT 28.600 30.200 28.900 31.800 ;
        RECT 23.800 29.800 24.200 30.200 ;
        RECT 28.600 29.800 29.000 30.200 ;
        RECT 21.400 27.100 21.800 27.200 ;
        RECT 22.200 27.100 22.600 27.200 ;
        RECT 21.400 26.800 22.600 27.100 ;
        RECT 19.800 25.800 20.200 26.200 ;
        RECT 23.800 24.200 24.100 29.800 ;
        RECT 35.000 27.200 35.300 36.800 ;
        RECT 37.400 34.800 37.800 35.200 ;
        RECT 44.600 34.800 45.000 35.200 ;
        RECT 47.800 34.800 48.200 35.200 ;
        RECT 37.400 34.200 37.700 34.800 ;
        RECT 37.400 33.800 37.800 34.200 ;
        RECT 36.600 32.800 37.000 33.200 ;
        RECT 27.000 26.800 27.400 27.200 ;
        RECT 29.400 27.100 29.800 27.200 ;
        RECT 30.200 27.100 30.600 27.200 ;
        RECT 29.400 26.800 30.600 27.100 ;
        RECT 35.000 26.800 35.400 27.200 ;
        RECT 27.000 24.200 27.300 26.800 ;
        RECT 36.600 26.200 36.900 32.800 ;
        RECT 44.600 30.200 44.900 34.800 ;
        RECT 47.800 34.200 48.100 34.800 ;
        RECT 47.000 33.800 47.400 34.200 ;
        RECT 47.800 33.800 48.200 34.200 ;
        RECT 45.400 31.800 45.800 32.200 ;
        RECT 44.600 29.800 45.000 30.200 ;
        RECT 38.200 28.800 38.600 29.200 ;
        RECT 40.600 28.800 41.000 29.200 ;
        RECT 38.200 26.200 38.500 28.800 ;
        RECT 39.000 27.800 39.400 28.200 ;
        RECT 39.000 27.200 39.300 27.800 ;
        RECT 39.000 26.800 39.400 27.200 ;
        RECT 36.600 25.800 37.000 26.200 ;
        RECT 38.200 25.800 38.600 26.200 ;
        RECT 34.200 24.800 34.600 25.200 ;
        RECT 34.200 24.200 34.500 24.800 ;
        RECT 40.600 24.200 40.900 28.800 ;
        RECT 44.600 26.200 44.900 29.800 ;
        RECT 45.400 29.200 45.700 31.800 ;
        RECT 45.400 28.800 45.800 29.200 ;
        RECT 47.000 27.200 47.300 33.800 ;
        RECT 46.200 26.800 46.600 27.200 ;
        RECT 47.000 26.800 47.400 27.200 ;
        RECT 46.200 26.200 46.500 26.800 ;
        RECT 42.200 25.800 42.600 26.200 ;
        RECT 44.600 25.800 45.000 26.200 ;
        RECT 46.200 25.800 46.600 26.200 ;
        RECT 42.200 25.200 42.500 25.800 ;
        RECT 42.200 24.800 42.600 25.200 ;
        RECT 43.000 24.800 43.400 25.200 ;
        RECT 43.000 24.200 43.300 24.800 ;
        RECT 19.000 24.100 19.400 24.200 ;
        RECT 19.800 24.100 20.200 24.200 ;
        RECT 19.000 23.800 20.200 24.100 ;
        RECT 23.800 23.800 24.200 24.200 ;
        RECT 25.400 23.800 25.800 24.200 ;
        RECT 27.000 23.800 27.400 24.200 ;
        RECT 34.200 23.800 34.600 24.200 ;
        RECT 40.600 23.800 41.000 24.200 ;
        RECT 43.000 23.800 43.400 24.200 ;
        RECT 44.600 23.800 45.000 24.200 ;
        RECT 24.600 21.800 25.000 22.200 ;
        RECT 2.200 18.800 2.600 19.200 ;
        RECT 8.600 18.800 9.000 19.200 ;
        RECT 18.200 18.800 18.600 19.200 ;
        RECT 19.800 18.800 20.200 19.200 ;
        RECT 19.800 18.200 20.100 18.800 ;
        RECT 24.600 18.200 24.900 21.800 ;
        RECT 1.400 17.800 1.800 18.200 ;
        RECT 15.000 17.800 15.400 18.200 ;
        RECT 19.800 17.800 20.200 18.200 ;
        RECT 24.600 17.800 25.000 18.200 ;
        RECT 1.400 17.200 1.700 17.800 ;
        RECT 15.000 17.200 15.300 17.800 ;
        RECT 1.400 16.800 1.800 17.200 ;
        RECT 4.600 16.800 5.000 17.200 ;
        RECT 6.200 16.800 6.600 17.200 ;
        RECT 15.000 16.800 15.400 17.200 ;
        RECT 16.600 16.800 17.000 17.200 ;
        RECT 20.600 16.800 21.000 17.200 ;
        RECT 24.600 16.800 25.000 17.200 ;
        RECT 2.200 15.800 2.600 16.200 ;
        RECT 3.000 15.800 3.400 16.200 ;
        RECT 3.800 15.800 4.200 16.200 ;
        RECT 2.200 15.200 2.500 15.800 ;
        RECT 2.200 14.800 2.600 15.200 ;
        RECT 3.000 9.200 3.300 15.800 ;
        RECT 3.800 15.200 4.100 15.800 ;
        RECT 3.800 14.800 4.200 15.200 ;
        RECT 4.600 13.200 4.900 16.800 ;
        RECT 6.200 16.200 6.500 16.800 ;
        RECT 16.600 16.200 16.900 16.800 ;
        RECT 6.200 15.800 6.600 16.200 ;
        RECT 7.000 16.100 7.400 16.200 ;
        RECT 7.000 15.800 8.100 16.100 ;
        RECT 5.400 15.100 5.800 15.200 ;
        RECT 6.200 15.100 6.600 15.200 ;
        RECT 5.400 14.800 6.600 15.100 ;
        RECT 6.200 13.800 6.600 14.200 ;
        RECT 4.600 12.800 5.000 13.200 ;
        RECT 3.000 8.800 3.400 9.200 ;
        RECT 5.400 8.800 5.800 9.200 ;
        RECT 1.300 7.500 1.700 7.900 ;
        RECT 3.000 7.800 3.400 8.200 ;
        RECT 2.200 7.500 4.300 7.800 ;
        RECT 4.600 7.500 5.000 7.900 ;
        RECT 1.300 5.100 1.600 7.500 ;
        RECT 2.200 7.400 2.600 7.500 ;
        RECT 3.900 7.400 4.300 7.500 ;
        RECT 4.700 7.100 5.000 7.500 ;
        RECT 2.600 6.800 5.000 7.100 ;
        RECT 5.400 7.200 5.700 8.800 ;
        RECT 6.200 8.200 6.500 13.800 ;
        RECT 7.800 9.200 8.100 15.800 ;
        RECT 10.200 15.800 10.600 16.200 ;
        RECT 13.400 16.100 13.800 16.200 ;
        RECT 14.200 16.100 14.600 16.200 ;
        RECT 13.400 15.800 14.600 16.100 ;
        RECT 16.600 15.800 17.000 16.200 ;
        RECT 18.200 15.800 18.600 16.200 ;
        RECT 19.000 15.800 19.400 16.200 ;
        RECT 9.400 13.800 9.800 14.200 ;
        RECT 9.400 12.200 9.700 13.800 ;
        RECT 10.200 13.200 10.500 15.800 ;
        RECT 12.600 15.100 13.000 15.200 ;
        RECT 13.400 15.100 13.800 15.200 ;
        RECT 12.600 14.800 13.800 15.100 ;
        RECT 11.800 13.800 12.200 14.200 ;
        RECT 15.800 13.800 16.200 14.200 ;
        RECT 11.800 13.200 12.100 13.800 ;
        RECT 10.200 12.800 10.600 13.200 ;
        RECT 11.800 12.800 12.200 13.200 ;
        RECT 9.400 11.800 9.800 12.200 ;
        RECT 10.200 10.200 10.500 12.800 ;
        RECT 12.600 11.800 13.000 12.200 ;
        RECT 10.200 9.800 10.600 10.200 ;
        RECT 12.600 9.200 12.900 11.800 ;
        RECT 7.800 8.800 8.200 9.200 ;
        RECT 11.800 8.800 12.200 9.200 ;
        RECT 12.600 8.800 13.000 9.200 ;
        RECT 6.200 7.800 6.600 8.200 ;
        RECT 7.100 7.800 7.500 7.900 ;
        RECT 6.200 7.200 6.500 7.800 ;
        RECT 7.100 7.500 9.900 7.800 ;
        RECT 10.200 7.500 10.600 7.900 ;
        RECT 5.400 6.800 5.800 7.200 ;
        RECT 6.200 6.800 6.600 7.200 ;
        RECT 2.600 6.700 3.000 6.800 ;
        RECT 4.700 5.100 5.000 6.800 ;
        RECT 1.300 4.700 1.700 5.100 ;
        RECT 4.600 4.700 5.000 5.100 ;
        RECT 7.100 5.100 7.400 7.500 ;
        RECT 7.800 7.400 8.200 7.500 ;
        RECT 9.500 7.400 9.900 7.500 ;
        RECT 10.300 7.100 10.600 7.500 ;
        RECT 7.800 6.800 10.600 7.100 ;
        RECT 11.800 7.200 12.100 8.800 ;
        RECT 11.800 6.800 12.200 7.200 ;
        RECT 7.800 6.100 8.100 6.800 ;
        RECT 7.700 5.700 8.100 6.100 ;
        RECT 10.300 5.100 10.600 6.800 ;
        RECT 15.800 6.200 16.100 13.800 ;
        RECT 16.600 8.200 16.900 15.800 ;
        RECT 18.200 15.200 18.500 15.800 ;
        RECT 17.400 14.800 17.800 15.200 ;
        RECT 18.200 14.800 18.600 15.200 ;
        RECT 17.400 11.200 17.700 14.800 ;
        RECT 19.000 14.200 19.300 15.800 ;
        RECT 19.000 13.800 19.400 14.200 ;
        RECT 19.000 12.200 19.300 13.800 ;
        RECT 19.000 11.800 19.400 12.200 ;
        RECT 17.400 10.800 17.800 11.200 ;
        RECT 16.600 7.800 17.000 8.200 ;
        RECT 17.400 7.200 17.700 10.800 ;
        RECT 20.600 9.200 20.900 16.800 ;
        RECT 21.400 15.800 21.800 16.200 ;
        RECT 23.000 15.800 23.400 16.200 ;
        RECT 21.400 15.200 21.700 15.800 ;
        RECT 23.000 15.200 23.300 15.800 ;
        RECT 21.400 14.800 21.800 15.200 ;
        RECT 23.000 14.800 23.400 15.200 ;
        RECT 23.800 14.800 24.200 15.200 ;
        RECT 23.800 13.200 24.100 14.800 ;
        RECT 24.600 14.200 24.900 16.800 ;
        RECT 24.600 13.800 25.000 14.200 ;
        RECT 23.800 12.800 24.200 13.200 ;
        RECT 23.800 11.800 24.200 12.200 ;
        RECT 23.000 9.800 23.400 10.200 ;
        RECT 18.200 8.800 18.600 9.200 ;
        RECT 20.600 8.800 21.000 9.200 ;
        RECT 18.200 7.200 18.500 8.800 ;
        RECT 19.000 7.500 19.400 7.900 ;
        RECT 19.700 7.500 21.800 7.800 ;
        RECT 22.300 7.500 22.700 7.900 ;
        RECT 17.400 6.800 17.800 7.200 ;
        RECT 18.200 6.800 18.600 7.200 ;
        RECT 19.000 7.100 19.300 7.500 ;
        RECT 19.700 7.400 20.100 7.500 ;
        RECT 21.400 7.400 21.800 7.500 ;
        RECT 19.000 6.800 21.400 7.100 ;
        RECT 15.000 6.100 15.400 6.200 ;
        RECT 15.800 6.100 16.200 6.200 ;
        RECT 15.000 5.800 16.200 6.100 ;
        RECT 7.100 4.700 7.500 5.100 ;
        RECT 10.200 4.700 10.600 5.100 ;
        RECT 19.000 5.100 19.300 6.800 ;
        RECT 21.000 6.700 21.400 6.800 ;
        RECT 22.400 5.100 22.700 7.500 ;
        RECT 23.000 7.200 23.300 9.800 ;
        RECT 23.800 8.200 24.100 11.800 ;
        RECT 24.600 9.200 24.900 13.800 ;
        RECT 25.400 9.200 25.700 23.800 ;
        RECT 27.800 21.800 28.200 22.200 ;
        RECT 36.600 22.100 37.000 22.200 ;
        RECT 37.400 22.100 37.800 22.200 ;
        RECT 36.600 21.800 37.800 22.100 ;
        RECT 39.800 21.800 40.200 22.200 ;
        RECT 43.800 21.800 44.200 22.200 ;
        RECT 27.800 16.200 28.100 21.800 ;
        RECT 31.000 17.800 31.400 18.200 ;
        RECT 32.600 17.800 33.000 18.200 ;
        RECT 34.200 17.800 34.600 18.200 ;
        RECT 31.000 16.200 31.300 17.800 ;
        RECT 27.800 15.800 28.200 16.200 ;
        RECT 31.000 15.800 31.400 16.200 ;
        RECT 31.800 15.800 32.200 16.200 ;
        RECT 28.600 15.100 29.000 15.200 ;
        RECT 29.400 15.100 29.800 15.200 ;
        RECT 28.600 14.800 29.800 15.100 ;
        RECT 31.800 14.200 32.100 15.800 ;
        RECT 32.600 15.200 32.900 17.800 ;
        RECT 34.200 17.200 34.500 17.800 ;
        RECT 39.800 17.200 40.100 21.800 ;
        RECT 34.200 16.800 34.600 17.200 ;
        RECT 35.800 17.100 36.200 17.200 ;
        RECT 36.600 17.100 37.000 17.200 ;
        RECT 35.800 16.800 37.000 17.100 ;
        RECT 39.800 16.800 40.200 17.200 ;
        RECT 35.000 15.800 35.400 16.200 ;
        RECT 36.600 15.800 37.000 16.200 ;
        RECT 37.400 15.800 37.800 16.200 ;
        RECT 35.000 15.200 35.300 15.800 ;
        RECT 36.600 15.200 36.900 15.800 ;
        RECT 32.600 14.800 33.000 15.200 ;
        RECT 35.000 14.800 35.400 15.200 ;
        RECT 36.600 14.800 37.000 15.200 ;
        RECT 26.200 13.800 26.600 14.200 ;
        RECT 27.800 13.800 28.200 14.200 ;
        RECT 29.400 14.100 29.800 14.200 ;
        RECT 30.200 14.100 30.600 14.200 ;
        RECT 29.400 13.800 30.600 14.100 ;
        RECT 31.800 13.800 32.200 14.200 ;
        RECT 37.400 14.100 37.700 15.800 ;
        RECT 39.800 14.200 40.100 16.800 ;
        RECT 43.800 16.200 44.100 21.800 ;
        RECT 44.600 17.200 44.900 23.800 ;
        RECT 51.000 23.200 51.300 45.800 ;
        RECT 52.600 45.200 52.900 45.800 ;
        RECT 52.600 44.800 53.000 45.200 ;
        RECT 52.600 43.200 52.900 44.800 ;
        RECT 55.000 43.200 55.300 46.800 ;
        RECT 55.800 45.200 56.100 46.800 ;
        RECT 55.800 44.800 56.200 45.200 ;
        RECT 58.200 44.800 58.600 45.200 ;
        RECT 52.600 42.800 53.000 43.200 ;
        RECT 55.000 42.800 55.400 43.200 ;
        RECT 51.800 39.800 52.200 40.200 ;
        RECT 51.800 29.200 52.100 39.800 ;
        RECT 55.000 34.200 55.300 42.800 ;
        RECT 55.800 39.200 56.100 44.800 ;
        RECT 58.200 41.200 58.500 44.800 ;
        RECT 58.200 40.800 58.600 41.200 ;
        RECT 55.800 38.800 56.200 39.200 ;
        RECT 57.400 37.800 57.800 38.200 ;
        RECT 57.400 37.200 57.700 37.800 ;
        RECT 57.400 36.800 57.800 37.200 ;
        RECT 59.000 35.200 59.300 46.800 ;
        RECT 59.800 45.800 60.200 46.200 ;
        RECT 59.800 40.200 60.100 45.800 ;
        RECT 62.200 41.800 62.600 42.200 ;
        RECT 62.200 41.200 62.500 41.800 ;
        RECT 62.200 40.800 62.600 41.200 ;
        RECT 59.800 39.800 60.200 40.200 ;
        RECT 61.400 39.800 61.800 40.200 ;
        RECT 59.800 37.200 60.100 39.800 ;
        RECT 61.400 39.200 61.700 39.800 ;
        RECT 61.400 38.800 61.800 39.200 ;
        RECT 59.800 36.800 60.200 37.200 ;
        RECT 59.000 34.800 59.400 35.200 ;
        RECT 59.800 34.800 60.200 35.200 ;
        RECT 55.000 33.800 55.400 34.200 ;
        RECT 59.000 29.200 59.300 34.800 ;
        RECT 51.800 28.800 52.200 29.200 ;
        RECT 59.000 28.800 59.400 29.200 ;
        RECT 53.400 26.800 53.800 27.200 ;
        RECT 56.600 26.800 57.000 27.200 ;
        RECT 58.200 27.100 58.600 27.200 ;
        RECT 59.800 27.100 60.100 34.800 ;
        RECT 62.200 29.800 62.600 30.200 ;
        RECT 62.200 28.200 62.500 29.800 ;
        RECT 63.000 29.200 63.300 49.800 ;
        RECT 63.800 47.200 64.100 51.800 ;
        RECT 64.600 49.200 64.900 54.800 ;
        RECT 64.600 48.800 65.000 49.200 ;
        RECT 65.400 48.200 65.700 66.800 ;
        RECT 67.000 65.800 67.400 66.200 ;
        RECT 67.000 56.200 67.300 65.800 ;
        RECT 71.800 64.800 72.200 65.200 ;
        RECT 68.600 63.800 69.000 64.200 ;
        RECT 67.000 55.800 67.400 56.200 ;
        RECT 67.000 55.200 67.300 55.800 ;
        RECT 68.600 55.200 68.900 63.800 ;
        RECT 71.800 58.200 72.100 64.800 ;
        RECT 72.600 63.200 72.900 73.800 ;
        RECT 73.400 69.200 73.700 80.800 ;
        RECT 75.000 79.800 75.400 80.200 ;
        RECT 77.400 79.800 77.800 80.200 ;
        RECT 74.200 77.800 74.600 78.200 ;
        RECT 74.200 76.200 74.500 77.800 ;
        RECT 74.200 75.800 74.600 76.200 ;
        RECT 75.000 75.200 75.300 79.800 ;
        RECT 77.400 79.200 77.700 79.800 ;
        RECT 77.400 78.800 77.800 79.200 ;
        RECT 80.600 78.200 80.900 86.800 ;
        RECT 81.400 86.100 81.800 86.200 ;
        RECT 82.200 86.100 82.600 86.200 ;
        RECT 81.400 85.800 82.600 86.100 ;
        RECT 87.000 85.200 87.300 87.800 ;
        RECT 88.600 86.800 89.000 87.200 ;
        RECT 89.400 86.800 89.800 87.200 ;
        RECT 91.000 87.100 91.400 87.200 ;
        RECT 91.800 87.100 92.200 87.200 ;
        RECT 91.000 86.800 92.200 87.100 ;
        RECT 93.400 86.800 93.800 87.200 ;
        RECT 87.000 84.800 87.400 85.200 ;
        RECT 87.000 82.800 87.400 83.200 ;
        RECT 83.800 82.100 84.200 82.200 ;
        RECT 84.600 82.100 85.000 82.200 ;
        RECT 83.800 81.800 85.000 82.100 ;
        RECT 81.400 79.800 81.800 80.200 ;
        RECT 80.600 77.800 81.000 78.200 ;
        RECT 75.800 77.100 76.200 77.200 ;
        RECT 76.600 77.100 77.000 77.200 ;
        RECT 75.800 76.800 77.000 77.100 ;
        RECT 75.000 74.800 75.400 75.200 ;
        RECT 80.600 74.800 81.000 75.200 ;
        RECT 75.000 74.200 75.300 74.800 ;
        RECT 80.600 74.200 80.900 74.800 ;
        RECT 81.400 74.200 81.700 79.800 ;
        RECT 82.200 78.800 82.600 79.200 ;
        RECT 82.200 78.200 82.500 78.800 ;
        RECT 82.200 77.800 82.600 78.200 ;
        RECT 84.600 75.800 85.000 76.200 ;
        RECT 85.400 76.100 85.800 76.200 ;
        RECT 86.200 76.100 86.600 76.200 ;
        RECT 85.400 75.800 86.600 76.100 ;
        RECT 75.000 73.800 75.400 74.200 ;
        RECT 76.600 73.800 77.000 74.200 ;
        RECT 80.600 73.800 81.000 74.200 ;
        RECT 81.400 73.800 81.800 74.200 ;
        RECT 83.000 73.800 83.400 74.200 ;
        RECT 83.800 73.800 84.200 74.200 ;
        RECT 73.400 68.800 73.800 69.200 ;
        RECT 75.000 68.800 75.400 69.200 ;
        RECT 75.000 67.200 75.300 68.800 ;
        RECT 75.000 66.800 75.400 67.200 ;
        RECT 74.200 65.800 74.600 66.200 ;
        RECT 75.000 65.800 75.400 66.200 ;
        RECT 76.600 66.100 76.900 73.800 ;
        RECT 81.400 73.200 81.700 73.800 ;
        RECT 81.400 72.800 81.800 73.200 ;
        RECT 83.000 72.200 83.300 73.800 ;
        RECT 83.800 73.200 84.100 73.800 ;
        RECT 83.800 72.800 84.200 73.200 ;
        RECT 78.200 71.800 78.600 72.200 ;
        RECT 79.800 71.800 80.200 72.200 ;
        RECT 83.000 71.800 83.400 72.200 ;
        RECT 78.200 66.200 78.500 71.800 ;
        RECT 77.400 66.100 77.800 66.200 ;
        RECT 76.600 65.800 77.800 66.100 ;
        RECT 78.200 65.800 78.600 66.200 ;
        RECT 72.600 62.800 73.000 63.200 ;
        RECT 71.800 57.800 72.200 58.200 ;
        RECT 67.000 54.800 67.400 55.200 ;
        RECT 68.600 54.800 69.000 55.200 ;
        RECT 72.600 55.100 73.000 55.200 ;
        RECT 73.400 55.100 73.800 55.200 ;
        RECT 72.600 54.800 73.800 55.100 ;
        RECT 67.000 53.800 67.400 54.200 ;
        RECT 67.000 53.200 67.300 53.800 ;
        RECT 67.000 52.800 67.400 53.200 ;
        RECT 67.800 51.800 68.200 52.200 ;
        RECT 67.800 49.200 68.100 51.800 ;
        RECT 67.800 48.800 68.200 49.200 ;
        RECT 65.400 47.800 65.800 48.200 ;
        RECT 63.800 46.800 64.200 47.200 ;
        RECT 68.600 44.200 68.900 54.800 ;
        RECT 71.000 53.800 71.400 54.200 ;
        RECT 71.000 53.200 71.300 53.800 ;
        RECT 69.400 52.800 69.800 53.200 ;
        RECT 71.000 52.800 71.400 53.200 ;
        RECT 69.400 49.200 69.700 52.800 ;
        RECT 70.200 50.800 70.600 51.200 ;
        RECT 71.800 50.800 72.200 51.200 ;
        RECT 70.200 49.200 70.500 50.800 ;
        RECT 69.400 48.800 69.800 49.200 ;
        RECT 70.200 48.800 70.600 49.200 ;
        RECT 69.400 48.200 69.700 48.800 ;
        RECT 69.400 47.800 69.800 48.200 ;
        RECT 71.800 47.200 72.100 50.800 ;
        RECT 72.600 47.800 73.000 48.200 ;
        RECT 72.600 47.200 72.900 47.800 ;
        RECT 74.200 47.200 74.500 65.800 ;
        RECT 75.000 61.200 75.300 65.800 ;
        RECT 76.600 63.200 76.900 65.800 ;
        RECT 77.400 65.100 77.800 65.200 ;
        RECT 78.200 65.100 78.500 65.800 ;
        RECT 77.400 64.800 78.500 65.100 ;
        RECT 76.600 62.800 77.000 63.200 ;
        RECT 76.600 62.200 76.900 62.800 ;
        RECT 79.800 62.200 80.100 71.800 ;
        RECT 84.600 69.200 84.900 75.800 ;
        RECT 86.200 74.800 86.600 75.200 ;
        RECT 86.200 72.200 86.500 74.800 ;
        RECT 87.000 74.200 87.300 82.800 ;
        RECT 87.800 81.800 88.200 82.200 ;
        RECT 87.800 79.200 88.100 81.800 ;
        RECT 87.800 78.800 88.200 79.200 ;
        RECT 88.600 77.200 88.900 86.800 ;
        RECT 89.400 86.200 89.700 86.800 ;
        RECT 89.400 85.800 89.800 86.200 ;
        RECT 91.000 84.800 91.400 85.200 ;
        RECT 91.000 83.200 91.300 84.800 ;
        RECT 93.400 83.200 93.700 86.800 ;
        RECT 91.000 82.800 91.400 83.200 ;
        RECT 93.400 82.800 93.800 83.200 ;
        RECT 94.200 78.200 94.500 87.800 ;
        RECT 96.600 86.200 96.900 93.800 ;
        RECT 96.600 85.800 97.000 86.200 ;
        RECT 96.600 82.200 96.900 85.800 ;
        RECT 95.800 81.800 96.200 82.200 ;
        RECT 96.600 81.800 97.000 82.200 ;
        RECT 89.400 77.800 89.800 78.200 ;
        RECT 94.200 77.800 94.600 78.200 ;
        RECT 88.600 76.800 89.000 77.200 ;
        RECT 89.400 74.200 89.700 77.800 ;
        RECT 91.800 76.800 92.200 77.200 ;
        RECT 91.800 76.200 92.100 76.800 ;
        RECT 94.200 76.200 94.500 77.800 ;
        RECT 95.800 77.200 96.100 81.800 ;
        RECT 95.800 76.800 96.200 77.200 ;
        RECT 91.800 75.800 92.200 76.200 ;
        RECT 94.200 75.800 94.600 76.200 ;
        RECT 95.000 75.800 95.400 76.200 ;
        RECT 90.200 74.800 90.600 75.200 ;
        RECT 90.200 74.200 90.500 74.800 ;
        RECT 95.000 74.200 95.300 75.800 ;
        RECT 95.800 74.800 96.200 75.200 ;
        RECT 87.000 73.800 87.400 74.200 ;
        RECT 89.400 73.800 89.800 74.200 ;
        RECT 90.200 73.800 90.600 74.200 ;
        RECT 92.600 73.800 93.000 74.200 ;
        RECT 94.200 73.800 94.600 74.200 ;
        RECT 95.000 73.800 95.400 74.200 ;
        RECT 88.600 72.800 89.000 73.200 ;
        RECT 91.800 72.800 92.200 73.200 ;
        RECT 86.200 71.800 86.600 72.200 ;
        RECT 87.000 70.800 87.400 71.200 ;
        RECT 87.000 69.200 87.300 70.800 ;
        RECT 84.600 68.800 85.000 69.200 ;
        RECT 87.000 68.800 87.400 69.200 ;
        RECT 88.600 65.200 88.900 72.800 ;
        RECT 91.800 72.200 92.100 72.800 ;
        RECT 91.800 71.800 92.200 72.200 ;
        RECT 92.600 66.200 92.900 73.800 ;
        RECT 94.200 73.200 94.500 73.800 ;
        RECT 94.200 72.800 94.600 73.200 ;
        RECT 95.800 73.100 96.100 74.800 ;
        RECT 95.000 72.800 96.100 73.100 ;
        RECT 95.000 72.200 95.300 72.800 ;
        RECT 95.000 71.800 95.400 72.200 ;
        RECT 95.800 71.800 96.200 72.200 ;
        RECT 95.800 69.200 96.100 71.800 ;
        RECT 95.800 68.800 96.200 69.200 ;
        RECT 96.600 68.100 96.900 81.800 ;
        RECT 97.400 76.200 97.700 95.800 ;
        RECT 99.000 94.800 99.400 95.200 ;
        RECT 98.200 93.800 98.600 94.200 ;
        RECT 98.200 92.200 98.500 93.800 ;
        RECT 99.000 93.200 99.300 94.800 ;
        RECT 99.000 92.800 99.400 93.200 ;
        RECT 98.200 91.800 98.600 92.200 ;
        RECT 97.400 75.800 97.800 76.200 ;
        RECT 98.200 71.200 98.500 91.800 ;
        RECT 102.200 89.200 102.500 95.800 ;
        RECT 103.800 94.800 104.200 95.200 ;
        RECT 105.400 94.800 105.800 95.200 ;
        RECT 107.000 95.100 107.400 95.200 ;
        RECT 107.800 95.100 108.200 95.200 ;
        RECT 107.000 94.800 108.200 95.100 ;
        RECT 110.200 94.800 110.600 95.200 ;
        RECT 115.800 94.800 116.200 95.200 ;
        RECT 118.200 94.800 118.600 95.200 ;
        RECT 103.800 94.200 104.100 94.800 ;
        RECT 105.400 94.200 105.700 94.800 ;
        RECT 103.000 93.800 103.400 94.200 ;
        RECT 103.800 93.800 104.200 94.200 ;
        RECT 105.400 93.800 105.800 94.200 ;
        RECT 103.000 93.200 103.300 93.800 ;
        RECT 103.000 92.800 103.400 93.200 ;
        RECT 102.200 88.800 102.600 89.200 ;
        RECT 106.200 88.800 106.600 89.200 ;
        RECT 106.200 88.200 106.500 88.800 ;
        RECT 101.400 87.500 101.800 87.900 ;
        RECT 102.100 87.500 104.200 87.800 ;
        RECT 104.700 87.500 105.100 87.900 ;
        RECT 106.200 87.800 106.600 88.200 ;
        RECT 101.400 87.100 101.700 87.500 ;
        RECT 102.100 87.400 102.500 87.500 ;
        RECT 103.800 87.400 104.200 87.500 ;
        RECT 101.400 86.800 103.800 87.100 ;
        RECT 101.400 85.100 101.700 86.800 ;
        RECT 103.400 86.700 103.800 86.800 ;
        RECT 101.400 84.700 101.800 85.100 ;
        RECT 103.800 84.800 104.200 85.200 ;
        RECT 104.800 85.100 105.100 87.500 ;
        RECT 105.400 87.100 105.800 87.200 ;
        RECT 106.200 87.100 106.600 87.200 ;
        RECT 105.400 86.800 106.600 87.100 ;
        RECT 103.800 79.200 104.100 84.800 ;
        RECT 104.700 84.700 105.100 85.100 ;
        RECT 107.000 79.200 107.300 94.800 ;
        RECT 110.200 94.200 110.500 94.800 ;
        RECT 110.200 93.800 110.600 94.200 ;
        RECT 114.200 93.800 114.600 94.200 ;
        RECT 114.200 93.200 114.500 93.800 ;
        RECT 109.400 92.800 109.800 93.200 ;
        RECT 111.800 93.100 112.200 93.200 ;
        RECT 111.800 92.800 112.900 93.100 ;
        RECT 114.200 92.800 114.600 93.200 ;
        RECT 109.400 92.200 109.700 92.800 ;
        RECT 109.400 91.800 109.800 92.200 ;
        RECT 109.400 90.200 109.700 91.800 ;
        RECT 109.400 89.800 109.800 90.200 ;
        RECT 112.600 89.200 112.900 92.800 ;
        RECT 115.800 92.200 116.100 94.800 ;
        RECT 118.200 94.200 118.500 94.800 ;
        RECT 118.200 93.800 118.600 94.200 ;
        RECT 119.000 94.100 119.400 94.200 ;
        RECT 119.800 94.100 120.200 94.200 ;
        RECT 119.000 93.800 120.200 94.100 ;
        RECT 121.400 93.200 121.700 101.800 ;
        RECT 122.200 94.200 122.500 114.800 ;
        RECT 124.600 114.800 125.000 115.200 ;
        RECT 123.000 107.100 123.400 107.200 ;
        RECT 123.800 107.100 124.200 107.200 ;
        RECT 123.000 106.800 124.200 107.100 ;
        RECT 124.600 106.200 124.900 114.800 ;
        RECT 126.200 112.100 126.600 118.900 ;
        RECT 127.000 112.100 127.400 118.900 ;
        RECT 127.800 112.100 128.200 117.900 ;
        RECT 128.600 115.800 129.000 116.200 ;
        RECT 128.600 114.200 128.900 115.800 ;
        RECT 128.600 113.800 129.000 114.200 ;
        RECT 129.400 112.100 129.800 117.900 ;
        RECT 131.000 112.100 131.400 117.900 ;
        RECT 131.800 112.100 132.200 118.900 ;
        RECT 132.600 112.100 133.000 118.900 ;
        RECT 133.400 112.100 133.800 118.900 ;
        RECT 140.600 115.200 140.900 120.800 ;
        RECT 140.600 114.800 141.000 115.200 ;
        RECT 143.800 114.800 144.200 115.200 ;
        RECT 146.200 114.800 146.600 115.200 ;
        RECT 139.000 114.100 139.400 114.200 ;
        RECT 139.800 114.100 140.200 114.200 ;
        RECT 139.000 113.800 140.200 114.100 ;
        RECT 140.600 113.800 141.000 114.200 ;
        RECT 140.600 113.200 140.900 113.800 ;
        RECT 143.800 113.200 144.100 114.800 ;
        RECT 139.800 112.800 140.200 113.200 ;
        RECT 140.600 113.100 141.000 113.200 ;
        RECT 141.400 113.100 141.800 113.200 ;
        RECT 140.600 112.800 141.800 113.100 ;
        RECT 143.800 112.800 144.200 113.200 ;
        RECT 139.800 112.200 140.100 112.800 ;
        RECT 139.800 111.800 140.200 112.200 ;
        RECT 124.600 105.800 125.000 106.200 ;
        RECT 127.000 105.800 127.400 106.200 ;
        RECT 124.600 104.200 124.900 105.800 ;
        RECT 124.600 103.800 125.000 104.200 ;
        RECT 127.000 95.200 127.300 105.800 ;
        RECT 127.800 102.100 128.200 108.900 ;
        RECT 128.600 102.100 129.000 108.900 ;
        RECT 129.400 103.100 129.800 108.900 ;
        RECT 130.200 107.800 130.600 108.200 ;
        RECT 130.200 107.200 130.500 107.800 ;
        RECT 130.200 106.800 130.600 107.200 ;
        RECT 131.000 103.100 131.400 108.900 ;
        RECT 132.600 103.100 133.000 108.900 ;
        RECT 133.400 102.100 133.800 108.900 ;
        RECT 134.200 102.100 134.600 108.900 ;
        RECT 135.000 102.100 135.400 108.900 ;
        RECT 139.800 105.200 140.100 111.800 ;
        RECT 145.400 109.800 145.800 110.200 ;
        RECT 145.400 108.100 145.700 109.800 ;
        RECT 146.200 109.100 146.500 114.800 ;
        RECT 147.000 111.200 147.300 121.800 ;
        RECT 147.000 110.800 147.400 111.200 ;
        RECT 147.000 109.100 147.400 109.200 ;
        RECT 146.200 108.800 147.400 109.100 ;
        RECT 146.200 108.100 146.600 108.200 ;
        RECT 145.400 107.800 146.600 108.100 ;
        RECT 141.400 106.800 141.800 107.200 ;
        RECT 146.200 106.800 146.600 107.200 ;
        RECT 141.400 106.200 141.700 106.800 ;
        RECT 146.200 106.200 146.500 106.800 ;
        RECT 141.400 106.100 141.800 106.200 ;
        RECT 142.200 106.100 142.600 106.200 ;
        RECT 141.400 105.800 142.600 106.100 ;
        RECT 143.000 106.100 143.400 106.200 ;
        RECT 143.800 106.100 144.200 106.200 ;
        RECT 143.000 105.800 144.200 106.100 ;
        RECT 146.200 105.800 146.600 106.200 ;
        RECT 147.000 106.100 147.400 106.200 ;
        RECT 147.800 106.100 148.200 106.200 ;
        RECT 147.000 105.800 148.200 106.100 ;
        RECT 139.800 104.800 140.200 105.200 ;
        RECT 142.200 105.100 142.600 105.200 ;
        RECT 143.000 105.100 143.400 105.200 ;
        RECT 142.200 104.800 143.400 105.100 ;
        RECT 140.600 103.800 141.000 104.200 ;
        RECT 144.600 103.800 145.000 104.200 ;
        RECT 127.000 94.800 127.400 95.200 ;
        RECT 122.200 93.800 122.600 94.200 ;
        RECT 121.400 93.100 121.800 93.200 ;
        RECT 122.200 93.100 122.600 93.200 ;
        RECT 121.400 92.800 122.600 93.100 ;
        RECT 115.800 91.800 116.200 92.200 ;
        RECT 124.600 91.800 125.000 92.200 ;
        RECT 127.800 92.100 128.200 98.900 ;
        RECT 128.600 92.100 129.000 98.900 ;
        RECT 129.400 92.100 129.800 97.900 ;
        RECT 130.200 93.800 130.600 94.200 ;
        RECT 124.600 89.200 124.900 91.800 ;
        RECT 128.600 89.800 129.000 90.200 ;
        RECT 112.600 88.800 113.000 89.200 ;
        RECT 119.800 88.800 120.200 89.200 ;
        RECT 124.600 88.800 125.000 89.200 ;
        RECT 119.800 88.200 120.100 88.800 ;
        RECT 117.400 88.100 117.800 88.200 ;
        RECT 118.200 88.100 118.600 88.200 ;
        RECT 117.400 87.800 118.600 88.100 ;
        RECT 119.000 87.800 119.400 88.200 ;
        RECT 119.800 87.800 120.200 88.200 ;
        RECT 123.800 87.800 124.200 88.200 ;
        RECT 124.600 87.800 125.000 88.200 ;
        RECT 125.400 87.800 125.800 88.200 ;
        RECT 126.200 87.800 126.600 88.200 ;
        RECT 107.800 86.800 108.200 87.200 ;
        RECT 109.400 87.100 109.800 87.200 ;
        RECT 110.200 87.100 110.600 87.200 ;
        RECT 109.400 86.800 110.600 87.100 ;
        RECT 111.000 86.800 111.400 87.200 ;
        RECT 111.800 86.800 112.200 87.200 ;
        RECT 115.800 87.100 116.200 87.200 ;
        RECT 116.600 87.100 117.000 87.200 ;
        RECT 115.800 86.800 117.000 87.100 ;
        RECT 107.800 80.200 108.100 86.800 ;
        RECT 111.000 86.200 111.300 86.800 ;
        RECT 111.000 85.800 111.400 86.200 ;
        RECT 111.800 84.100 112.100 86.800 ;
        RECT 119.000 86.200 119.300 87.800 ;
        RECT 123.800 87.200 124.100 87.800 ;
        RECT 120.600 86.800 121.000 87.200 ;
        RECT 122.200 87.100 122.600 87.200 ;
        RECT 123.000 87.100 123.400 87.200 ;
        RECT 122.200 86.800 123.400 87.100 ;
        RECT 123.800 86.800 124.200 87.200 ;
        RECT 116.600 86.100 117.000 86.200 ;
        RECT 117.400 86.100 117.800 86.200 ;
        RECT 116.600 85.800 117.800 86.100 ;
        RECT 119.000 85.800 119.400 86.200 ;
        RECT 111.000 83.800 112.100 84.100 ;
        RECT 114.200 84.800 114.600 85.200 ;
        RECT 114.200 84.200 114.500 84.800 ;
        RECT 114.200 83.800 114.600 84.200 ;
        RECT 108.600 82.100 109.000 82.200 ;
        RECT 109.400 82.100 109.800 82.200 ;
        RECT 108.600 81.800 109.800 82.100 ;
        RECT 107.800 79.800 108.200 80.200 ;
        RECT 111.000 79.200 111.300 83.800 ;
        RECT 112.600 80.800 113.000 81.200 ;
        RECT 102.200 78.800 102.600 79.200 ;
        RECT 103.800 78.800 104.200 79.200 ;
        RECT 107.000 78.800 107.400 79.200 ;
        RECT 111.000 78.800 111.400 79.200 ;
        RECT 99.000 74.800 99.400 75.200 ;
        RECT 101.400 74.800 101.800 75.200 ;
        RECT 99.000 74.200 99.300 74.800 ;
        RECT 99.000 73.800 99.400 74.200 ;
        RECT 101.400 73.200 101.700 74.800 ;
        RECT 101.400 72.800 101.800 73.200 ;
        RECT 99.000 71.800 99.400 72.200 ;
        RECT 98.200 70.800 98.600 71.200 ;
        RECT 99.000 69.100 99.300 71.800 ;
        RECT 99.000 68.800 100.100 69.100 ;
        RECT 95.800 67.800 96.900 68.100 ;
        RECT 98.200 67.800 98.600 68.200 ;
        RECT 99.000 67.800 99.400 68.200 ;
        RECT 94.200 66.800 94.600 67.200 ;
        RECT 91.000 66.100 91.400 66.200 ;
        RECT 91.800 66.100 92.200 66.200 ;
        RECT 91.000 65.800 92.200 66.100 ;
        RECT 92.600 65.800 93.000 66.200 ;
        RECT 84.600 64.800 85.000 65.200 ;
        RECT 87.000 65.100 87.400 65.200 ;
        RECT 86.200 64.800 87.400 65.100 ;
        RECT 88.600 64.800 89.000 65.200 ;
        RECT 90.200 64.800 90.600 65.200 ;
        RECT 75.800 61.800 76.200 62.200 ;
        RECT 76.600 61.800 77.000 62.200 ;
        RECT 79.800 61.800 80.200 62.200 ;
        RECT 80.600 61.800 81.000 62.200 ;
        RECT 75.000 60.800 75.400 61.200 ;
        RECT 75.000 56.200 75.300 60.800 ;
        RECT 75.800 56.200 76.100 61.800 ;
        RECT 80.600 58.200 80.900 61.800 ;
        RECT 84.600 60.200 84.900 64.800 ;
        RECT 84.600 59.800 85.000 60.200 ;
        RECT 79.000 57.800 79.400 58.200 ;
        RECT 80.600 57.800 81.000 58.200 ;
        RECT 79.000 57.200 79.300 57.800 ;
        RECT 79.000 56.800 79.400 57.200 ;
        RECT 75.000 55.800 75.400 56.200 ;
        RECT 75.800 55.800 76.200 56.200 ;
        RECT 77.400 55.800 77.800 56.200 ;
        RECT 80.600 56.100 81.000 56.200 ;
        RECT 81.400 56.100 81.800 56.200 ;
        RECT 80.600 55.800 81.800 56.100 ;
        RECT 75.000 53.200 75.300 55.800 ;
        RECT 75.000 52.800 75.400 53.200 ;
        RECT 75.800 52.100 76.200 52.200 ;
        RECT 76.600 52.100 77.000 52.200 ;
        RECT 75.800 51.800 77.000 52.100 ;
        RECT 77.400 49.200 77.700 55.800 ;
        RECT 86.200 55.200 86.500 64.800 ;
        RECT 90.200 64.200 90.500 64.800 ;
        RECT 90.200 63.800 90.600 64.200 ;
        RECT 92.600 63.200 92.900 65.800 ;
        RECT 94.200 65.200 94.500 66.800 ;
        RECT 94.200 64.800 94.600 65.200 ;
        RECT 92.600 62.800 93.000 63.200 ;
        RECT 92.600 62.100 93.000 62.200 ;
        RECT 93.400 62.100 93.800 62.200 ;
        RECT 92.600 61.800 93.800 62.100 ;
        RECT 91.000 59.800 91.400 60.200 ;
        RECT 87.000 56.100 87.400 56.200 ;
        RECT 87.800 56.100 88.200 56.200 ;
        RECT 87.000 55.800 88.200 56.100 ;
        RECT 79.000 54.800 79.400 55.200 ;
        RECT 79.800 54.800 80.200 55.200 ;
        RECT 83.000 54.800 83.400 55.200 ;
        RECT 86.200 54.800 86.600 55.200 ;
        RECT 79.000 51.200 79.300 54.800 ;
        RECT 79.800 54.200 80.100 54.800 ;
        RECT 79.800 53.800 80.200 54.200 ;
        RECT 79.000 50.800 79.400 51.200 ;
        RECT 77.400 48.800 77.800 49.200 ;
        RECT 82.200 48.800 82.600 49.200 ;
        RECT 75.000 47.800 75.400 48.200 ;
        RECT 79.800 47.800 80.200 48.200 ;
        RECT 69.400 47.100 69.800 47.200 ;
        RECT 70.200 47.100 70.600 47.200 ;
        RECT 69.400 46.800 70.600 47.100 ;
        RECT 71.000 47.100 71.400 47.200 ;
        RECT 71.800 47.100 72.200 47.200 ;
        RECT 71.000 46.800 72.200 47.100 ;
        RECT 72.600 46.800 73.000 47.200 ;
        RECT 74.200 47.100 74.600 47.200 ;
        RECT 75.000 47.100 75.300 47.800 ;
        RECT 74.200 46.800 75.300 47.100 ;
        RECT 74.200 44.800 74.600 45.200 ;
        RECT 68.600 43.800 69.000 44.200 ;
        RECT 68.600 41.800 69.000 42.200 ;
        RECT 71.000 41.800 71.400 42.200 ;
        RECT 73.400 41.800 73.800 42.200 ;
        RECT 68.600 35.200 68.900 41.800 ;
        RECT 71.000 36.200 71.300 41.800 ;
        RECT 71.800 38.800 72.200 39.200 ;
        RECT 71.000 35.800 71.400 36.200 ;
        RECT 71.800 35.200 72.100 38.800 ;
        RECT 73.400 36.200 73.700 41.800 ;
        RECT 74.200 39.200 74.500 44.800 ;
        RECT 74.200 38.800 74.600 39.200 ;
        RECT 73.400 35.800 73.800 36.200 ;
        RECT 75.000 35.200 75.300 46.800 ;
        RECT 77.400 46.800 77.800 47.200 ;
        RECT 79.000 46.800 79.400 47.200 ;
        RECT 75.800 46.100 76.200 46.200 ;
        RECT 76.600 46.100 77.000 46.200 ;
        RECT 75.800 45.800 77.000 46.100 ;
        RECT 75.800 44.800 76.200 45.200 ;
        RECT 75.800 39.200 76.100 44.800 ;
        RECT 77.400 42.200 77.700 46.800 ;
        RECT 79.000 46.200 79.300 46.800 ;
        RECT 78.200 45.800 78.600 46.200 ;
        RECT 79.000 45.800 79.400 46.200 ;
        RECT 78.200 45.200 78.500 45.800 ;
        RECT 78.200 44.800 78.600 45.200 ;
        RECT 76.600 41.800 77.000 42.200 ;
        RECT 77.400 41.800 77.800 42.200 ;
        RECT 76.600 40.200 76.900 41.800 ;
        RECT 77.400 40.800 77.800 41.200 ;
        RECT 76.600 39.800 77.000 40.200 ;
        RECT 75.800 38.800 76.200 39.200 ;
        RECT 77.400 37.200 77.700 40.800 ;
        RECT 79.800 39.200 80.100 47.800 ;
        RECT 82.200 47.200 82.500 48.800 ;
        RECT 80.600 47.100 81.000 47.200 ;
        RECT 81.400 47.100 81.800 47.200 ;
        RECT 80.600 46.800 81.800 47.100 ;
        RECT 82.200 46.800 82.600 47.200 ;
        RECT 83.000 46.200 83.300 54.800 ;
        RECT 85.400 53.800 85.800 54.200 ;
        RECT 85.400 52.200 85.700 53.800 ;
        RECT 83.800 51.800 84.200 52.200 ;
        RECT 85.400 51.800 85.800 52.200 ;
        RECT 83.800 51.200 84.100 51.800 ;
        RECT 83.800 50.800 84.200 51.200 ;
        RECT 86.200 48.200 86.500 54.800 ;
        RECT 87.800 53.200 88.100 55.800 ;
        RECT 91.000 55.200 91.300 59.800 ;
        RECT 92.600 56.800 93.000 57.200 ;
        RECT 92.600 56.200 92.900 56.800 ;
        RECT 95.800 56.200 96.100 67.800 ;
        RECT 98.200 67.200 98.500 67.800 ;
        RECT 96.600 66.800 97.000 67.200 ;
        RECT 98.200 66.800 98.600 67.200 ;
        RECT 96.600 66.200 96.900 66.800 ;
        RECT 96.600 65.800 97.000 66.200 ;
        RECT 99.000 65.200 99.300 67.800 ;
        RECT 99.000 64.800 99.400 65.200 ;
        RECT 92.600 55.800 93.000 56.200 ;
        RECT 95.800 55.800 96.200 56.200 ;
        RECT 98.200 55.800 98.600 56.200 ;
        RECT 88.600 54.800 89.000 55.200 ;
        RECT 91.000 54.800 91.400 55.200 ;
        RECT 93.400 55.100 93.800 55.200 ;
        RECT 94.200 55.100 94.600 55.200 ;
        RECT 93.400 54.800 94.600 55.100 ;
        RECT 88.600 54.200 88.900 54.800 ;
        RECT 88.600 53.800 89.000 54.200 ;
        RECT 89.400 54.100 89.800 54.200 ;
        RECT 90.200 54.100 90.600 54.200 ;
        RECT 89.400 53.800 90.600 54.100 ;
        RECT 93.400 53.800 93.800 54.200 ;
        RECT 95.000 53.800 95.400 54.200 ;
        RECT 93.400 53.200 93.700 53.800 ;
        RECT 87.800 52.800 88.200 53.200 ;
        RECT 93.400 52.800 93.800 53.200 ;
        RECT 89.400 51.800 89.800 52.200 ;
        RECT 92.600 51.800 93.000 52.200 ;
        RECT 86.200 47.800 86.600 48.200 ;
        RECT 87.800 47.800 88.200 48.200 ;
        RECT 89.400 48.100 89.700 51.800 ;
        RECT 92.600 48.200 92.900 51.800 ;
        RECT 89.400 47.800 90.500 48.100 ;
        RECT 92.600 47.800 93.000 48.200 ;
        RECT 87.800 47.200 88.100 47.800 ;
        RECT 90.200 47.200 90.500 47.800 ;
        RECT 83.800 46.800 84.200 47.200 ;
        RECT 87.800 46.800 88.200 47.200 ;
        RECT 88.600 47.100 89.000 47.200 ;
        RECT 89.400 47.100 89.800 47.200 ;
        RECT 88.600 46.800 89.800 47.100 ;
        RECT 90.200 46.800 90.600 47.200 ;
        RECT 92.600 47.100 93.000 47.200 ;
        RECT 93.400 47.100 93.800 47.200 ;
        RECT 92.600 46.800 93.800 47.100 ;
        RECT 81.400 45.800 81.800 46.200 ;
        RECT 83.000 45.800 83.400 46.200 ;
        RECT 81.400 44.200 81.700 45.800 ;
        RECT 83.000 44.800 83.400 45.200 ;
        RECT 81.400 43.800 81.800 44.200 ;
        RECT 81.400 43.200 81.700 43.800 ;
        RECT 81.400 42.800 81.800 43.200 ;
        RECT 79.800 38.800 80.200 39.200 ;
        RECT 77.400 36.800 77.800 37.200 ;
        RECT 80.600 36.800 81.000 37.200 ;
        RECT 68.600 35.100 69.000 35.200 ;
        RECT 69.400 35.100 69.800 35.200 ;
        RECT 68.600 34.800 69.800 35.100 ;
        RECT 70.200 35.100 70.600 35.200 ;
        RECT 71.000 35.100 71.400 35.200 ;
        RECT 70.200 34.800 71.400 35.100 ;
        RECT 71.800 34.800 72.200 35.200 ;
        RECT 75.000 35.100 75.400 35.200 ;
        RECT 75.800 35.100 76.200 35.200 ;
        RECT 75.000 34.800 76.200 35.100 ;
        RECT 79.800 34.800 80.200 35.200 ;
        RECT 69.400 34.200 69.700 34.800 ;
        RECT 79.800 34.200 80.100 34.800 ;
        RECT 80.600 34.200 80.900 36.800 ;
        RECT 82.200 35.800 82.600 36.200 ;
        RECT 82.200 35.200 82.500 35.800 ;
        RECT 83.000 35.200 83.300 44.800 ;
        RECT 83.800 37.200 84.100 46.800 ;
        RECT 95.000 46.200 95.300 53.800 ;
        RECT 95.800 50.200 96.100 55.800 ;
        RECT 98.200 55.200 98.500 55.800 ;
        RECT 96.600 55.100 97.000 55.200 ;
        RECT 97.400 55.100 97.800 55.200 ;
        RECT 96.600 54.800 97.800 55.100 ;
        RECT 98.200 54.800 98.600 55.200 ;
        RECT 95.800 49.800 96.200 50.200 ;
        RECT 97.400 49.800 97.800 50.200 ;
        RECT 95.800 46.800 96.200 47.200 ;
        RECT 84.600 45.800 85.000 46.200 ;
        RECT 85.400 45.800 85.800 46.200 ;
        RECT 86.200 45.800 86.600 46.200 ;
        RECT 88.600 45.800 89.000 46.200 ;
        RECT 91.000 46.100 91.400 46.200 ;
        RECT 91.800 46.100 92.200 46.200 ;
        RECT 91.000 45.800 92.200 46.100 ;
        RECT 95.000 45.800 95.400 46.200 ;
        RECT 84.600 38.200 84.900 45.800 ;
        RECT 85.400 45.200 85.700 45.800 ;
        RECT 86.200 45.200 86.500 45.800 ;
        RECT 85.400 44.800 85.800 45.200 ;
        RECT 86.200 44.800 86.600 45.200 ;
        RECT 87.000 44.800 87.400 45.200 ;
        RECT 87.000 43.200 87.300 44.800 ;
        RECT 85.400 42.800 85.800 43.200 ;
        RECT 87.000 42.800 87.400 43.200 ;
        RECT 85.400 39.200 85.700 42.800 ;
        RECT 88.600 42.200 88.900 45.800 ;
        RECT 95.000 45.200 95.300 45.800 ;
        RECT 95.800 45.200 96.100 46.800 ;
        RECT 97.400 46.200 97.700 49.800 ;
        RECT 99.000 49.200 99.300 64.800 ;
        RECT 99.800 63.200 100.100 68.800 ;
        RECT 101.400 66.800 101.800 67.200 ;
        RECT 99.800 62.800 100.200 63.200 ;
        RECT 101.400 60.200 101.700 66.800 ;
        RECT 102.200 66.200 102.500 78.800 ;
        RECT 107.800 76.800 108.200 77.200 ;
        RECT 107.800 75.200 108.100 76.800 ;
        RECT 105.400 74.800 105.800 75.200 ;
        RECT 107.800 74.800 108.200 75.200 ;
        RECT 103.000 73.800 103.400 74.200 ;
        RECT 103.000 71.200 103.300 73.800 ;
        RECT 105.400 73.200 105.700 74.800 ;
        RECT 107.000 73.800 107.400 74.200 ;
        RECT 108.600 73.800 109.000 74.200 ;
        RECT 104.600 72.800 105.000 73.200 ;
        RECT 105.400 72.800 105.800 73.200 ;
        RECT 103.000 70.800 103.400 71.200 ;
        RECT 104.600 68.100 104.900 72.800 ;
        RECT 105.400 71.800 105.800 72.200 ;
        RECT 106.200 71.800 106.600 72.200 ;
        RECT 105.400 69.200 105.700 71.800 ;
        RECT 105.400 68.800 105.800 69.200 ;
        RECT 104.600 67.800 105.700 68.100 ;
        RECT 103.800 67.100 104.200 67.200 ;
        RECT 104.600 67.100 105.000 67.200 ;
        RECT 103.800 66.800 105.000 67.100 ;
        RECT 102.200 65.800 102.600 66.200 ;
        RECT 104.600 65.800 105.000 66.200 ;
        RECT 104.600 65.200 104.900 65.800 ;
        RECT 103.800 64.800 104.200 65.200 ;
        RECT 104.600 64.800 105.000 65.200 ;
        RECT 101.400 59.800 101.800 60.200 ;
        RECT 100.600 57.800 101.000 58.200 ;
        RECT 100.600 54.200 100.900 57.800 ;
        RECT 101.400 56.800 101.800 57.200 ;
        RECT 101.400 56.200 101.700 56.800 ;
        RECT 101.400 55.800 101.800 56.200 ;
        RECT 101.400 54.800 101.800 55.200 ;
        RECT 101.400 54.200 101.700 54.800 ;
        RECT 103.800 54.200 104.100 64.800 ;
        RECT 105.400 58.200 105.700 67.800 ;
        RECT 106.200 67.100 106.500 71.800 ;
        RECT 107.000 71.200 107.300 73.800 ;
        RECT 107.000 70.800 107.400 71.200 ;
        RECT 106.200 66.800 107.300 67.100 ;
        RECT 106.200 65.800 106.600 66.200 ;
        RECT 106.200 65.200 106.500 65.800 ;
        RECT 107.000 65.200 107.300 66.800 ;
        RECT 108.600 66.200 108.900 73.800 ;
        RECT 111.000 73.100 111.400 73.200 ;
        RECT 111.800 73.100 112.200 73.200 ;
        RECT 111.000 72.800 112.200 73.100 ;
        RECT 111.800 72.200 112.100 72.800 ;
        RECT 110.200 71.800 110.600 72.200 ;
        RECT 111.800 71.800 112.200 72.200 ;
        RECT 109.400 67.100 109.800 67.200 ;
        RECT 110.200 67.100 110.500 71.800 ;
        RECT 109.400 66.800 110.500 67.100 ;
        RECT 111.000 70.800 111.400 71.200 ;
        RECT 108.600 65.800 109.000 66.200 ;
        RECT 106.200 64.800 106.600 65.200 ;
        RECT 107.000 64.800 107.400 65.200 ;
        RECT 110.200 65.100 110.600 65.200 ;
        RECT 111.000 65.100 111.300 70.800 ;
        RECT 111.800 67.800 112.200 68.200 ;
        RECT 111.800 66.200 112.100 67.800 ;
        RECT 112.600 67.200 112.900 80.800 ;
        RECT 119.000 79.800 119.400 80.200 ;
        RECT 119.000 79.200 119.300 79.800 ;
        RECT 119.000 78.800 119.400 79.200 ;
        RECT 120.600 77.200 120.900 86.800 ;
        RECT 123.000 85.800 123.400 86.200 ;
        RECT 122.200 78.800 122.600 79.200 ;
        RECT 120.600 76.800 121.000 77.200 ;
        RECT 121.400 76.800 121.800 77.200 ;
        RECT 121.400 76.200 121.700 76.800 ;
        RECT 114.200 75.800 114.600 76.200 ;
        RECT 121.400 75.800 121.800 76.200 ;
        RECT 113.400 74.800 113.800 75.200 ;
        RECT 113.400 74.200 113.700 74.800 ;
        RECT 114.200 74.200 114.500 75.800 ;
        RECT 115.000 74.800 115.400 75.200 ;
        RECT 119.000 74.800 119.400 75.200 ;
        RECT 119.800 74.800 120.200 75.200 ;
        RECT 113.400 73.800 113.800 74.200 ;
        RECT 114.200 73.800 114.600 74.200 ;
        RECT 115.000 73.200 115.300 74.800 ;
        RECT 119.000 74.200 119.300 74.800 ;
        RECT 119.000 73.800 119.400 74.200 ;
        RECT 115.000 72.800 115.400 73.200 ;
        RECT 116.600 72.800 117.000 73.200 ;
        RECT 116.600 70.200 116.900 72.800 ;
        RECT 119.800 72.200 120.100 74.800 ;
        RECT 122.200 74.200 122.500 78.800 ;
        RECT 123.000 74.200 123.300 85.800 ;
        RECT 123.800 81.800 124.200 82.200 ;
        RECT 121.400 73.800 121.800 74.200 ;
        RECT 122.200 73.800 122.600 74.200 ;
        RECT 123.000 73.800 123.400 74.200 ;
        RECT 120.600 72.800 121.000 73.200 ;
        RECT 119.800 71.800 120.200 72.200 ;
        RECT 115.000 70.100 115.400 70.200 ;
        RECT 114.200 69.800 115.400 70.100 ;
        RECT 116.600 69.800 117.000 70.200 ;
        RECT 114.200 69.200 114.500 69.800 ;
        RECT 114.200 68.800 114.600 69.200 ;
        RECT 115.000 68.100 115.400 68.200 ;
        RECT 115.800 68.100 116.200 68.200 ;
        RECT 115.000 67.800 116.200 68.100 ;
        RECT 117.400 67.800 117.800 68.200 ;
        RECT 118.200 67.800 118.600 68.200 ;
        RECT 119.000 67.800 119.400 68.200 ;
        RECT 117.400 67.200 117.700 67.800 ;
        RECT 112.600 66.800 113.000 67.200 ;
        RECT 115.000 66.800 115.400 67.200 ;
        RECT 117.400 66.800 117.800 67.200 ;
        RECT 111.800 65.800 112.200 66.200 ;
        RECT 112.600 65.800 113.000 66.200 ;
        RECT 110.200 64.800 111.300 65.100 ;
        RECT 112.600 65.200 112.900 65.800 ;
        RECT 112.600 64.800 113.000 65.200 ;
        RECT 105.400 57.800 105.800 58.200 ;
        RECT 105.400 55.200 105.700 57.800 ;
        RECT 106.200 55.200 106.500 64.800 ;
        RECT 108.600 61.800 109.000 62.200 ;
        RECT 108.600 56.200 108.900 61.800 ;
        RECT 111.800 60.800 112.200 61.200 ;
        RECT 111.000 56.800 111.400 57.200 ;
        RECT 108.600 55.800 109.000 56.200 ;
        RECT 110.200 55.800 110.600 56.200 ;
        RECT 110.200 55.200 110.500 55.800 ;
        RECT 105.400 54.800 105.800 55.200 ;
        RECT 106.200 54.800 106.600 55.200 ;
        RECT 107.000 54.800 107.400 55.200 ;
        RECT 110.200 54.800 110.600 55.200 ;
        RECT 100.600 53.800 101.000 54.200 ;
        RECT 101.400 53.800 101.800 54.200 ;
        RECT 103.800 53.800 104.200 54.200 ;
        RECT 104.600 54.100 105.000 54.200 ;
        RECT 105.400 54.100 105.800 54.200 ;
        RECT 104.600 53.800 105.800 54.100 ;
        RECT 103.000 53.100 103.400 53.200 ;
        RECT 103.800 53.100 104.200 53.200 ;
        RECT 103.000 52.800 104.200 53.100 ;
        RECT 104.600 52.800 105.000 53.200 ;
        RECT 105.400 52.800 105.800 53.200 ;
        RECT 107.000 53.100 107.300 54.800 ;
        RECT 111.000 54.200 111.300 56.800 ;
        RECT 111.800 55.200 112.100 60.800 ;
        RECT 115.000 57.200 115.300 66.800 ;
        RECT 115.800 66.100 116.200 66.200 ;
        RECT 116.600 66.100 117.000 66.200 ;
        RECT 115.800 65.800 117.000 66.100 ;
        RECT 118.200 65.200 118.500 67.800 ;
        RECT 119.000 66.200 119.300 67.800 ;
        RECT 120.600 67.200 120.900 72.800 ;
        RECT 121.400 67.200 121.700 73.800 ;
        RECT 122.200 73.100 122.600 73.200 ;
        RECT 123.000 73.100 123.400 73.200 ;
        RECT 122.200 72.800 123.400 73.100 ;
        RECT 123.800 72.200 124.100 81.800 ;
        RECT 124.600 74.200 124.900 87.800 ;
        RECT 125.400 87.200 125.700 87.800 ;
        RECT 126.200 87.200 126.500 87.800 ;
        RECT 125.400 86.800 125.800 87.200 ;
        RECT 126.200 86.800 126.600 87.200 ;
        RECT 127.800 86.800 128.200 87.200 ;
        RECT 127.800 86.200 128.100 86.800 ;
        RECT 128.600 86.200 128.900 89.800 ;
        RECT 130.200 89.200 130.500 93.800 ;
        RECT 131.000 92.100 131.400 97.900 ;
        RECT 132.600 92.100 133.000 97.900 ;
        RECT 133.400 92.100 133.800 98.900 ;
        RECT 134.200 92.100 134.600 98.900 ;
        RECT 135.000 92.100 135.400 98.900 ;
        RECT 139.900 95.800 140.300 96.200 ;
        RECT 139.900 95.200 140.200 95.800 ;
        RECT 140.600 95.200 140.900 103.800 ;
        RECT 144.600 99.200 144.900 103.800 ;
        RECT 144.600 98.800 145.000 99.200 ;
        RECT 148.600 95.200 148.900 121.800 ;
        RECT 139.900 94.800 140.300 95.200 ;
        RECT 140.600 94.800 141.000 95.200 ;
        RECT 143.800 94.800 144.200 95.200 ;
        RECT 145.400 94.800 145.800 95.200 ;
        RECT 146.200 95.100 146.600 95.200 ;
        RECT 147.000 95.100 147.400 95.200 ;
        RECT 146.200 94.800 147.400 95.100 ;
        RECT 148.600 94.800 149.000 95.200 ;
        RECT 139.800 93.800 140.200 94.200 ;
        RECT 139.800 89.200 140.100 93.800 ;
        RECT 143.800 93.200 144.100 94.800 ;
        RECT 145.400 94.100 145.700 94.800 ;
        RECT 145.400 93.800 146.500 94.100 ;
        RECT 145.400 93.200 145.700 93.800 ;
        RECT 143.800 92.800 144.200 93.200 ;
        RECT 145.400 92.800 145.800 93.200 ;
        RECT 130.200 88.800 130.600 89.200 ;
        RECT 139.800 88.800 140.200 89.200 ;
        RECT 140.600 89.100 141.000 89.200 ;
        RECT 141.400 89.100 141.800 89.200 ;
        RECT 140.600 88.800 141.800 89.100 ;
        RECT 143.800 88.200 144.100 92.800 ;
        RECT 131.000 87.800 131.400 88.200 ;
        RECT 131.000 87.200 131.300 87.800 ;
        RECT 133.300 87.500 133.700 87.900 ;
        RECT 134.200 87.500 136.300 87.800 ;
        RECT 136.600 87.500 137.000 87.900 ;
        RECT 129.400 86.800 129.800 87.200 ;
        RECT 131.000 86.800 131.400 87.200 ;
        RECT 131.800 87.100 132.200 87.200 ;
        RECT 132.600 87.100 133.000 87.200 ;
        RECT 131.800 86.800 133.000 87.100 ;
        RECT 126.200 86.100 126.600 86.200 ;
        RECT 127.000 86.100 127.400 86.200 ;
        RECT 126.200 85.800 127.400 86.100 ;
        RECT 127.800 85.800 128.200 86.200 ;
        RECT 128.600 85.800 129.000 86.200 ;
        RECT 128.600 84.800 129.000 85.200 ;
        RECT 128.600 83.200 128.900 84.800 ;
        RECT 128.600 82.800 129.000 83.200 ;
        RECT 127.000 78.800 127.400 79.200 ;
        RECT 127.000 75.200 127.300 78.800 ;
        RECT 128.600 77.800 129.000 78.200 ;
        RECT 128.600 77.200 128.900 77.800 ;
        RECT 128.600 76.800 129.000 77.200 ;
        RECT 129.400 76.200 129.700 86.800 ;
        RECT 130.200 85.800 130.600 86.200 ;
        RECT 130.200 76.200 130.500 85.800 ;
        RECT 131.800 84.800 132.200 85.200 ;
        RECT 133.300 85.100 133.600 87.500 ;
        RECT 134.200 87.400 134.600 87.500 ;
        RECT 135.900 87.400 136.300 87.500 ;
        RECT 136.700 87.100 137.000 87.500 ;
        RECT 140.600 87.800 141.000 88.200 ;
        RECT 143.800 87.800 144.200 88.200 ;
        RECT 144.600 88.100 145.000 88.200 ;
        RECT 145.400 88.100 145.800 88.200 ;
        RECT 144.600 87.800 145.800 88.100 ;
        RECT 134.600 86.800 137.000 87.100 ;
        RECT 134.600 86.700 135.000 86.800 ;
        RECT 135.800 85.800 136.200 86.200 ;
        RECT 135.800 85.200 136.100 85.800 ;
        RECT 131.800 79.200 132.100 84.800 ;
        RECT 133.300 84.700 133.700 85.100 ;
        RECT 135.800 84.800 136.200 85.200 ;
        RECT 136.700 85.100 137.000 86.800 ;
        RECT 136.600 84.700 137.000 85.100 ;
        RECT 137.400 86.800 137.800 87.200 ;
        RECT 139.000 86.800 139.400 87.200 ;
        RECT 137.400 85.200 137.700 86.800 ;
        RECT 139.000 86.200 139.300 86.800 ;
        RECT 138.200 85.800 138.600 86.200 ;
        RECT 139.000 85.800 139.400 86.200 ;
        RECT 137.400 84.800 137.800 85.200 ;
        RECT 138.200 84.200 138.500 85.800 ;
        RECT 138.200 83.800 138.600 84.200 ;
        RECT 135.800 79.800 136.200 80.200 ;
        RECT 131.000 78.800 131.400 79.200 ;
        RECT 131.800 78.800 132.200 79.200 ;
        RECT 129.400 75.800 129.800 76.200 ;
        RECT 130.200 75.800 130.600 76.200 ;
        RECT 129.400 75.200 129.700 75.800 ;
        RECT 125.400 74.800 125.800 75.200 ;
        RECT 127.000 74.800 127.400 75.200 ;
        RECT 129.400 74.800 129.800 75.200 ;
        RECT 125.400 74.200 125.700 74.800 ;
        RECT 124.600 73.800 125.000 74.200 ;
        RECT 125.400 73.800 125.800 74.200 ;
        RECT 126.200 73.800 126.600 74.200 ;
        RECT 129.400 74.100 129.800 74.200 ;
        RECT 130.200 74.100 130.600 74.200 ;
        RECT 129.400 73.800 130.600 74.100 ;
        RECT 126.200 72.200 126.500 73.800 ;
        RECT 123.800 71.800 124.200 72.200 ;
        RECT 126.200 71.800 126.600 72.200 ;
        RECT 123.800 68.200 124.100 71.800 ;
        RECT 130.200 70.800 130.600 71.200 ;
        RECT 130.200 69.200 130.500 70.800 ;
        RECT 128.600 68.800 129.000 69.200 ;
        RECT 130.200 68.800 130.600 69.200 ;
        RECT 122.200 68.100 122.600 68.200 ;
        RECT 123.000 68.100 123.400 68.200 ;
        RECT 122.200 67.800 123.400 68.100 ;
        RECT 123.800 67.800 124.200 68.200 ;
        RECT 126.200 67.800 126.600 68.200 ;
        RECT 127.000 67.800 127.400 68.200 ;
        RECT 126.200 67.200 126.500 67.800 ;
        RECT 127.000 67.200 127.300 67.800 ;
        RECT 128.600 67.200 128.900 68.800 ;
        RECT 131.000 68.200 131.300 78.800 ;
        RECT 132.600 76.800 133.000 77.200 ;
        RECT 134.200 76.800 134.600 77.200 ;
        RECT 132.600 76.200 132.900 76.800 ;
        RECT 131.800 75.800 132.200 76.200 ;
        RECT 132.600 75.800 133.000 76.200 ;
        RECT 131.800 74.200 132.100 75.800 ;
        RECT 134.200 75.200 134.500 76.800 ;
        RECT 135.800 76.200 136.100 79.800 ;
        RECT 136.600 77.800 137.000 78.200 ;
        RECT 137.400 77.800 137.800 78.200 ;
        RECT 135.800 75.800 136.200 76.200 ;
        RECT 134.200 74.800 134.600 75.200 ;
        RECT 135.800 74.800 136.200 75.200 ;
        RECT 135.800 74.200 136.100 74.800 ;
        RECT 136.600 74.200 136.900 77.800 ;
        RECT 137.400 77.200 137.700 77.800 ;
        RECT 137.400 76.800 137.800 77.200 ;
        RECT 137.400 75.800 137.800 76.200 ;
        RECT 139.000 75.800 139.400 76.200 ;
        RECT 137.400 75.200 137.700 75.800 ;
        RECT 139.000 75.200 139.300 75.800 ;
        RECT 137.400 74.800 137.800 75.200 ;
        RECT 139.000 74.800 139.400 75.200 ;
        RECT 131.800 73.800 132.200 74.200 ;
        RECT 132.600 74.100 133.000 74.200 ;
        RECT 133.400 74.100 133.800 74.200 ;
        RECT 132.600 73.800 133.800 74.100 ;
        RECT 135.800 73.800 136.200 74.200 ;
        RECT 136.600 73.800 137.000 74.200 ;
        RECT 133.400 68.800 133.800 69.200 ;
        RECT 131.000 67.800 131.400 68.200 ;
        RECT 131.800 67.800 132.200 68.200 ;
        RECT 131.800 67.200 132.100 67.800 ;
        RECT 133.400 67.200 133.700 68.800 ;
        RECT 136.600 68.100 136.900 73.800 ;
        RECT 140.600 70.200 140.900 87.800 ;
        RECT 146.200 86.200 146.500 93.800 ;
        RECT 148.600 92.800 149.000 93.200 ;
        RECT 146.200 85.800 146.600 86.200 ;
        RECT 148.600 85.200 148.900 92.800 ;
        RECT 149.400 91.800 149.800 92.200 ;
        RECT 141.400 84.800 141.800 85.200 ;
        RECT 148.600 84.800 149.000 85.200 ;
        RECT 141.400 79.200 141.700 84.800 ;
        RECT 146.200 83.800 146.600 84.200 ;
        RECT 146.200 79.200 146.500 83.800 ;
        RECT 148.600 82.200 148.900 84.800 ;
        RECT 149.400 83.100 149.700 91.800 ;
        RECT 150.200 86.800 150.600 87.200 ;
        RECT 150.200 84.200 150.500 86.800 ;
        RECT 150.200 83.800 150.600 84.200 ;
        RECT 149.400 82.800 150.500 83.100 ;
        RECT 148.600 81.800 149.000 82.200 ;
        RECT 149.400 81.800 149.800 82.200 ;
        RECT 141.400 78.800 141.800 79.200 ;
        RECT 146.200 78.800 146.600 79.200 ;
        RECT 145.400 75.800 145.800 76.200 ;
        RECT 145.400 75.200 145.700 75.800 ;
        RECT 141.400 74.800 141.800 75.200 ;
        RECT 142.200 74.800 142.600 75.200 ;
        RECT 145.400 74.800 145.800 75.200 ;
        RECT 141.400 73.200 141.700 74.800 ;
        RECT 142.200 74.200 142.500 74.800 ;
        RECT 142.200 73.800 142.600 74.200 ;
        RECT 143.000 74.100 143.400 74.200 ;
        RECT 143.800 74.100 144.200 74.200 ;
        RECT 143.000 73.800 144.200 74.100 ;
        RECT 147.000 73.800 147.400 74.200 ;
        RECT 141.400 72.800 141.800 73.200 ;
        RECT 143.000 72.800 143.400 73.200 ;
        RECT 140.600 69.800 141.000 70.200 ;
        RECT 143.000 69.200 143.300 72.800 ;
        RECT 146.200 71.800 146.600 72.200 ;
        RECT 143.800 69.800 144.200 70.200 ;
        RECT 143.800 69.200 144.100 69.800 ;
        RECT 146.200 69.200 146.500 71.800 ;
        RECT 147.000 71.200 147.300 73.800 ;
        RECT 148.600 71.800 149.000 72.200 ;
        RECT 147.000 70.800 147.400 71.200 ;
        RECT 143.000 68.800 143.400 69.200 ;
        RECT 143.800 68.800 144.200 69.200 ;
        RECT 146.200 68.800 146.600 69.200 ;
        RECT 136.600 67.800 137.700 68.100 ;
        RECT 137.400 67.200 137.700 67.800 ;
        RECT 139.000 67.800 139.400 68.200 ;
        RECT 147.000 67.800 147.400 68.200 ;
        RECT 139.000 67.200 139.300 67.800 ;
        RECT 120.600 66.800 121.000 67.200 ;
        RECT 121.400 66.800 121.800 67.200 ;
        RECT 123.000 67.100 123.400 67.200 ;
        RECT 123.800 67.100 124.200 67.200 ;
        RECT 123.000 66.800 124.200 67.100 ;
        RECT 125.400 66.800 125.800 67.200 ;
        RECT 126.200 66.800 126.600 67.200 ;
        RECT 127.000 66.800 127.400 67.200 ;
        RECT 128.600 66.800 129.000 67.200 ;
        RECT 131.800 66.800 132.200 67.200 ;
        RECT 132.600 66.800 133.000 67.200 ;
        RECT 133.400 66.800 133.800 67.200 ;
        RECT 135.000 66.800 135.400 67.200 ;
        RECT 136.600 66.800 137.000 67.200 ;
        RECT 137.400 66.800 137.800 67.200 ;
        RECT 139.000 66.800 139.400 67.200 ;
        RECT 145.400 66.800 145.800 67.200 ;
        RECT 120.600 66.200 120.900 66.800 ;
        RECT 125.400 66.200 125.700 66.800 ;
        RECT 119.000 65.800 119.400 66.200 ;
        RECT 120.600 65.800 121.000 66.200 ;
        RECT 125.400 65.800 125.800 66.200 ;
        RECT 127.000 66.100 127.400 66.200 ;
        RECT 127.800 66.100 128.200 66.200 ;
        RECT 127.000 65.800 128.200 66.100 ;
        RECT 116.600 64.800 117.000 65.200 ;
        RECT 118.200 64.800 118.600 65.200 ;
        RECT 123.000 64.800 123.400 65.200 ;
        RECT 123.800 65.100 124.200 65.200 ;
        RECT 124.600 65.100 125.000 65.200 ;
        RECT 123.800 64.800 125.000 65.100 ;
        RECT 116.600 59.200 116.900 64.800 ;
        RECT 123.000 62.200 123.300 64.800 ;
        RECT 125.400 64.200 125.700 65.800 ;
        RECT 128.600 65.200 128.900 66.800 ;
        RECT 132.600 66.200 132.900 66.800 ;
        RECT 135.000 66.200 135.300 66.800 ;
        RECT 136.600 66.200 136.900 66.800 ;
        RECT 130.200 65.800 130.600 66.200 ;
        RECT 132.600 65.800 133.000 66.200 ;
        RECT 134.200 65.800 134.600 66.200 ;
        RECT 135.000 65.800 135.400 66.200 ;
        RECT 135.800 65.800 136.200 66.200 ;
        RECT 136.600 65.800 137.000 66.200 ;
        RECT 139.800 65.800 140.200 66.200 ;
        RECT 141.400 65.800 141.800 66.200 ;
        RECT 130.200 65.200 130.500 65.800 ;
        RECT 127.800 64.800 128.200 65.200 ;
        RECT 128.600 64.800 129.000 65.200 ;
        RECT 130.200 64.800 130.600 65.200 ;
        RECT 125.400 63.800 125.800 64.200 ;
        RECT 120.600 61.800 121.000 62.200 ;
        RECT 123.000 61.800 123.400 62.200 ;
        RECT 116.600 58.800 117.000 59.200 ;
        RECT 113.400 56.800 113.800 57.200 ;
        RECT 115.000 56.800 115.400 57.200 ;
        RECT 113.400 56.200 113.700 56.800 ;
        RECT 120.600 56.200 120.900 61.800 ;
        RECT 124.600 57.800 125.000 58.200 ;
        RECT 113.400 55.800 113.800 56.200 ;
        RECT 118.200 56.100 118.600 56.200 ;
        RECT 119.000 56.100 119.400 56.200 ;
        RECT 118.200 55.800 119.400 56.100 ;
        RECT 120.600 55.800 121.000 56.200 ;
        RECT 122.200 55.800 122.600 56.200 ;
        RECT 122.200 55.200 122.500 55.800 ;
        RECT 111.800 54.800 112.200 55.200 ;
        RECT 115.800 55.100 116.200 55.200 ;
        RECT 116.600 55.100 117.000 55.200 ;
        RECT 115.800 54.800 117.000 55.100 ;
        RECT 120.600 55.100 121.000 55.200 ;
        RECT 121.400 55.100 121.800 55.200 ;
        RECT 120.600 54.800 121.800 55.100 ;
        RECT 122.200 54.800 122.600 55.200 ;
        RECT 123.000 55.100 123.400 55.200 ;
        RECT 123.800 55.100 124.200 55.200 ;
        RECT 123.000 54.800 124.200 55.100 ;
        RECT 124.600 54.200 124.900 57.800 ;
        RECT 127.800 55.200 128.100 64.800 ;
        RECT 132.600 64.200 132.900 65.800 ;
        RECT 132.600 63.800 133.000 64.200 ;
        RECT 132.600 57.800 133.000 58.200 ;
        RECT 130.200 56.800 130.600 57.200 ;
        RECT 130.200 56.200 130.500 56.800 ;
        RECT 130.200 55.800 130.600 56.200 ;
        RECT 132.600 55.200 132.900 57.800 ;
        RECT 133.400 55.800 133.800 56.200 ;
        RECT 133.400 55.200 133.700 55.800 ;
        RECT 134.200 55.200 134.500 65.800 ;
        RECT 135.800 65.100 136.100 65.800 ;
        RECT 135.800 64.800 136.900 65.100 ;
        RECT 135.800 61.800 136.200 62.200 ;
        RECT 135.800 59.200 136.100 61.800 ;
        RECT 135.800 58.800 136.200 59.200 ;
        RECT 135.000 57.800 135.400 58.200 ;
        RECT 135.000 57.200 135.300 57.800 ;
        RECT 135.000 56.800 135.400 57.200 ;
        RECT 127.800 54.800 128.200 55.200 ;
        RECT 132.600 54.800 133.000 55.200 ;
        RECT 133.400 54.800 133.800 55.200 ;
        RECT 134.200 54.800 134.600 55.200 ;
        RECT 136.600 54.200 136.900 64.800 ;
        RECT 137.400 64.800 137.800 65.200 ;
        RECT 137.400 64.200 137.700 64.800 ;
        RECT 137.400 63.800 137.800 64.200 ;
        RECT 139.000 54.800 139.400 55.200 ;
        RECT 108.600 54.100 109.000 54.200 ;
        RECT 109.400 54.100 109.800 54.200 ;
        RECT 108.600 53.800 109.800 54.100 ;
        RECT 111.000 53.800 111.400 54.200 ;
        RECT 115.800 53.800 116.200 54.200 ;
        RECT 119.000 53.800 119.400 54.200 ;
        RECT 124.600 53.800 125.000 54.200 ;
        RECT 126.200 54.100 126.600 54.200 ;
        RECT 127.000 54.100 127.400 54.200 ;
        RECT 126.200 53.800 127.400 54.100 ;
        RECT 131.800 53.800 132.200 54.200 ;
        RECT 136.600 54.100 137.000 54.200 ;
        RECT 137.400 54.100 137.800 54.200 ;
        RECT 136.600 53.800 137.800 54.100 ;
        RECT 107.800 53.100 108.200 53.200 ;
        RECT 107.000 52.800 108.200 53.100 ;
        RECT 109.400 52.800 109.800 53.200 ;
        RECT 104.600 49.200 104.900 52.800 ;
        RECT 105.400 49.200 105.700 52.800 ;
        RECT 107.800 52.200 108.100 52.800 ;
        RECT 107.800 51.800 108.200 52.200 ;
        RECT 108.600 51.800 109.000 52.200 ;
        RECT 99.000 48.800 99.400 49.200 ;
        RECT 104.600 48.800 105.000 49.200 ;
        RECT 105.400 48.800 105.800 49.200 ;
        RECT 99.000 47.800 101.700 48.100 ;
        RECT 99.000 47.200 99.300 47.800 ;
        RECT 101.400 47.200 101.700 47.800 ;
        RECT 103.800 47.800 104.200 48.200 ;
        RECT 103.800 47.200 104.100 47.800 ;
        RECT 99.000 46.800 99.400 47.200 ;
        RECT 99.800 47.100 100.200 47.200 ;
        RECT 100.600 47.100 101.000 47.200 ;
        RECT 99.800 46.800 101.000 47.100 ;
        RECT 101.400 46.800 101.800 47.200 ;
        RECT 103.800 46.800 104.200 47.200 ;
        RECT 97.400 45.800 97.800 46.200 ;
        RECT 99.000 45.800 99.400 46.200 ;
        RECT 99.800 45.800 100.200 46.200 ;
        RECT 101.400 45.800 101.800 46.200 ;
        RECT 102.200 46.100 102.600 46.200 ;
        RECT 103.000 46.100 103.400 46.200 ;
        RECT 102.200 45.800 103.400 46.100 ;
        RECT 93.400 45.100 93.800 45.200 ;
        RECT 94.200 45.100 94.600 45.200 ;
        RECT 93.400 44.800 94.600 45.100 ;
        RECT 95.000 44.800 95.400 45.200 ;
        RECT 95.800 44.800 96.200 45.200 ;
        RECT 96.600 42.800 97.000 43.200 ;
        RECT 88.600 41.800 89.000 42.200 ;
        RECT 85.400 38.800 85.800 39.200 ;
        RECT 86.200 38.800 86.600 39.200 ;
        RECT 91.800 38.800 92.200 39.200 ;
        RECT 84.600 37.800 85.000 38.200 ;
        RECT 83.800 36.800 84.200 37.200 ;
        RECT 83.800 35.800 84.200 36.200 ;
        RECT 84.600 35.800 85.000 36.200 ;
        RECT 83.800 35.200 84.100 35.800 ;
        RECT 84.600 35.200 84.900 35.800 ;
        RECT 81.400 34.800 81.800 35.200 ;
        RECT 82.200 34.800 82.600 35.200 ;
        RECT 83.000 34.800 83.400 35.200 ;
        RECT 83.800 34.800 84.200 35.200 ;
        RECT 84.600 34.800 85.000 35.200 ;
        RECT 81.400 34.200 81.700 34.800 ;
        RECT 86.200 34.200 86.500 38.800 ;
        RECT 87.800 37.100 88.200 37.200 ;
        RECT 88.600 37.100 89.000 37.200 ;
        RECT 87.800 36.800 89.000 37.100 ;
        RECT 87.000 35.800 87.400 36.200 ;
        RECT 90.200 35.800 90.600 36.200 ;
        RECT 68.600 33.800 69.000 34.200 ;
        RECT 69.400 33.800 69.800 34.200 ;
        RECT 71.800 33.800 72.200 34.200 ;
        RECT 75.000 33.800 75.400 34.200 ;
        RECT 79.800 33.800 80.200 34.200 ;
        RECT 80.600 33.800 81.000 34.200 ;
        RECT 81.400 33.800 81.800 34.200 ;
        RECT 82.200 33.800 82.600 34.200 ;
        RECT 83.000 33.800 83.400 34.200 ;
        RECT 86.200 33.800 86.600 34.200 ;
        RECT 65.400 33.100 65.800 33.200 ;
        RECT 66.200 33.100 66.600 33.200 ;
        RECT 65.400 32.800 66.600 33.100 ;
        RECT 64.600 29.800 65.000 30.200 ;
        RECT 63.000 28.800 63.400 29.200 ;
        RECT 64.600 28.200 64.900 29.800 ;
        RECT 65.400 28.800 65.800 29.200 ;
        RECT 62.200 27.800 62.600 28.200 ;
        RECT 64.600 27.800 65.000 28.200 ;
        RECT 65.400 27.200 65.700 28.800 ;
        RECT 68.600 28.200 68.900 33.800 ;
        RECT 71.800 33.200 72.100 33.800 ;
        RECT 75.000 33.200 75.300 33.800 ;
        RECT 71.800 32.800 72.200 33.200 ;
        RECT 74.200 32.800 74.600 33.200 ;
        RECT 75.000 32.800 75.400 33.200 ;
        RECT 74.200 32.200 74.500 32.800 ;
        RECT 74.200 31.800 74.600 32.200 ;
        RECT 78.200 31.800 78.600 32.200 ;
        RECT 78.200 31.200 78.500 31.800 ;
        RECT 75.000 30.800 75.400 31.200 ;
        RECT 78.200 30.800 78.600 31.200 ;
        RECT 69.400 28.800 69.800 29.200 ;
        RECT 71.000 28.800 71.400 29.200 ;
        RECT 73.400 29.100 73.800 29.200 ;
        RECT 74.200 29.100 74.600 29.200 ;
        RECT 73.400 28.800 74.600 29.100 ;
        RECT 67.800 27.800 68.200 28.200 ;
        RECT 68.600 27.800 69.000 28.200 ;
        RECT 58.200 26.800 60.100 27.100 ;
        RECT 53.400 24.200 53.700 26.800 ;
        RECT 56.600 26.200 56.900 26.800 ;
        RECT 56.600 25.800 57.000 26.200 ;
        RECT 58.200 25.800 58.600 26.200 ;
        RECT 59.000 25.800 59.400 26.200 ;
        RECT 55.000 25.100 55.400 25.200 ;
        RECT 55.800 25.100 56.200 25.200 ;
        RECT 55.000 24.800 56.200 25.100 ;
        RECT 53.400 23.800 53.800 24.200 ;
        RECT 58.200 23.200 58.500 25.800 ;
        RECT 59.000 25.200 59.300 25.800 ;
        RECT 59.000 24.800 59.400 25.200 ;
        RECT 51.000 22.800 51.400 23.200 ;
        RECT 58.200 22.800 58.600 23.200 ;
        RECT 44.600 16.800 45.000 17.200 ;
        RECT 40.600 15.800 41.000 16.200 ;
        RECT 43.800 15.800 44.200 16.200 ;
        RECT 48.600 15.800 49.000 16.200 ;
        RECT 40.600 15.200 40.900 15.800 ;
        RECT 48.600 15.200 48.900 15.800 ;
        RECT 51.000 15.200 51.300 22.800 ;
        RECT 56.600 21.800 57.000 22.200 ;
        RECT 53.400 16.800 53.800 17.200 ;
        RECT 55.800 16.800 56.200 17.200 ;
        RECT 40.600 14.800 41.000 15.200 ;
        RECT 48.600 14.800 49.000 15.200 ;
        RECT 51.000 14.800 51.400 15.200 ;
        RECT 51.000 14.200 51.300 14.800 ;
        RECT 38.200 14.100 38.600 14.200 ;
        RECT 37.400 13.800 38.600 14.100 ;
        RECT 39.800 13.800 40.200 14.200 ;
        RECT 40.600 14.100 41.000 14.200 ;
        RECT 41.400 14.100 41.800 14.200 ;
        RECT 40.600 13.800 41.800 14.100 ;
        RECT 45.400 14.100 45.800 14.200 ;
        RECT 46.200 14.100 46.600 14.200 ;
        RECT 45.400 13.800 46.600 14.100 ;
        RECT 51.000 13.800 51.400 14.200 ;
        RECT 26.200 13.200 26.500 13.800 ;
        RECT 27.800 13.200 28.100 13.800 ;
        RECT 38.200 13.200 38.500 13.800 ;
        RECT 53.400 13.200 53.700 16.800 ;
        RECT 55.800 16.200 56.100 16.800 ;
        RECT 55.800 15.800 56.200 16.200 ;
        RECT 26.200 12.800 26.600 13.200 ;
        RECT 27.800 12.800 28.200 13.200 ;
        RECT 38.200 12.800 38.600 13.200 ;
        RECT 41.400 12.800 41.800 13.200 ;
        RECT 46.200 12.800 46.600 13.200 ;
        RECT 49.400 12.800 49.800 13.200 ;
        RECT 53.400 12.800 53.800 13.200 ;
        RECT 27.000 11.800 27.400 12.200 ;
        RECT 30.200 11.800 30.600 12.200 ;
        RECT 39.000 11.800 39.400 12.200 ;
        RECT 24.600 8.800 25.000 9.200 ;
        RECT 25.400 8.800 25.800 9.200 ;
        RECT 23.800 7.800 24.200 8.200 ;
        RECT 23.000 6.800 23.400 7.200 ;
        RECT 27.000 6.200 27.300 11.800 ;
        RECT 30.200 10.200 30.500 11.800 ;
        RECT 39.000 11.200 39.300 11.800 ;
        RECT 35.800 10.800 36.200 11.200 ;
        RECT 39.000 10.800 39.400 11.200 ;
        RECT 28.600 9.800 29.000 10.200 ;
        RECT 30.200 9.800 30.600 10.200 ;
        RECT 35.000 9.800 35.400 10.200 ;
        RECT 27.800 7.800 28.200 8.200 ;
        RECT 27.800 7.200 28.100 7.800 ;
        RECT 28.600 7.200 28.900 9.800 ;
        RECT 33.400 8.800 33.800 9.200 ;
        RECT 29.500 7.800 29.900 7.900 ;
        RECT 29.500 7.500 32.300 7.800 ;
        RECT 32.600 7.500 33.000 7.900 ;
        RECT 27.800 6.800 28.200 7.200 ;
        RECT 28.600 6.800 29.000 7.200 ;
        RECT 27.000 5.800 27.400 6.200 ;
        RECT 19.000 4.700 19.400 5.100 ;
        RECT 22.300 4.700 22.700 5.100 ;
        RECT 25.400 5.100 25.800 5.200 ;
        RECT 26.200 5.100 26.600 5.200 ;
        RECT 25.400 4.800 26.600 5.100 ;
        RECT 29.500 5.100 29.800 7.500 ;
        RECT 30.200 7.400 30.600 7.500 ;
        RECT 31.900 7.400 32.300 7.500 ;
        RECT 32.700 7.100 33.000 7.500 ;
        RECT 30.200 6.800 33.000 7.100 ;
        RECT 33.400 7.200 33.700 8.800 ;
        RECT 35.000 8.200 35.300 9.800 ;
        RECT 35.000 7.800 35.400 8.200 ;
        RECT 35.800 7.200 36.100 10.800 ;
        RECT 37.400 7.800 37.800 8.200 ;
        RECT 37.400 7.200 37.700 7.800 ;
        RECT 41.400 7.200 41.700 12.800 ;
        RECT 46.200 12.200 46.500 12.800 ;
        RECT 46.200 11.800 46.600 12.200 ;
        RECT 47.000 11.800 47.400 12.200 ;
        RECT 47.000 7.200 47.300 11.800 ;
        RECT 49.400 9.200 49.700 12.800 ;
        RECT 52.600 11.800 53.000 12.200 ;
        RECT 49.400 8.800 49.800 9.200 ;
        RECT 33.400 6.800 33.800 7.200 ;
        RECT 35.800 6.800 36.200 7.200 ;
        RECT 37.400 6.800 37.800 7.200 ;
        RECT 41.400 6.800 41.800 7.200 ;
        RECT 44.600 7.100 45.000 7.200 ;
        RECT 45.400 7.100 45.800 7.200 ;
        RECT 44.600 6.800 45.800 7.100 ;
        RECT 47.000 6.800 47.400 7.200 ;
        RECT 49.400 6.800 49.800 7.200 ;
        RECT 30.200 6.100 30.500 6.800 ;
        RECT 30.100 5.700 30.500 6.100 ;
        RECT 30.200 5.100 30.600 5.200 ;
        RECT 31.000 5.100 31.400 5.200 ;
        RECT 32.700 5.100 33.000 6.800 ;
        RECT 49.400 6.200 49.700 6.800 ;
        RECT 52.600 6.200 52.900 11.800 ;
        RECT 53.400 11.200 53.700 12.800 ;
        RECT 53.400 10.800 53.800 11.200 ;
        RECT 56.600 7.200 56.900 21.800 ;
        RECT 59.800 19.200 60.100 26.800 ;
        RECT 61.400 26.800 61.800 27.200 ;
        RECT 65.400 26.800 65.800 27.200 ;
        RECT 59.800 18.800 60.200 19.200 ;
        RECT 61.400 15.200 61.700 26.800 ;
        RECT 67.800 26.200 68.100 27.800 ;
        RECT 69.400 27.200 69.700 28.800 ;
        RECT 71.000 28.200 71.300 28.800 ;
        RECT 70.200 27.800 70.600 28.200 ;
        RECT 71.000 27.800 71.400 28.200 ;
        RECT 68.600 26.800 69.000 27.200 ;
        RECT 69.400 26.800 69.800 27.200 ;
        RECT 66.200 26.100 66.600 26.200 ;
        RECT 67.000 26.100 67.400 26.200 ;
        RECT 66.200 25.800 67.400 26.100 ;
        RECT 67.800 25.800 68.200 26.200 ;
        RECT 68.600 25.200 68.900 26.800 ;
        RECT 63.000 25.100 63.400 25.200 ;
        RECT 63.800 25.100 64.200 25.200 ;
        RECT 65.400 25.100 65.800 25.200 ;
        RECT 63.000 24.800 64.200 25.100 ;
        RECT 64.600 24.800 65.800 25.100 ;
        RECT 68.600 24.800 69.000 25.200 ;
        RECT 63.800 15.800 64.200 16.200 ;
        RECT 63.800 15.200 64.100 15.800 ;
        RECT 61.400 14.800 61.800 15.200 ;
        RECT 63.800 14.800 64.200 15.200 ;
        RECT 58.200 9.800 58.600 10.200 ;
        RECT 58.200 9.200 58.500 9.800 ;
        RECT 61.400 9.200 61.700 14.800 ;
        RECT 63.800 12.800 64.200 13.200 ;
        RECT 63.800 9.200 64.100 12.800 ;
        RECT 64.600 11.200 64.900 24.800 ;
        RECT 65.400 23.800 65.800 24.200 ;
        RECT 65.400 13.200 65.700 23.800 ;
        RECT 67.800 15.800 68.200 16.200 ;
        RECT 67.800 15.200 68.100 15.800 ;
        RECT 70.200 15.200 70.500 27.800 ;
        RECT 75.000 26.200 75.300 30.800 ;
        RECT 77.400 28.800 77.800 29.200 ;
        RECT 78.200 28.800 78.600 29.200 ;
        RECT 79.000 29.100 79.400 29.200 ;
        RECT 79.800 29.100 80.200 29.200 ;
        RECT 79.000 28.800 80.200 29.100 ;
        RECT 75.800 26.800 76.200 27.200 ;
        RECT 77.400 27.100 77.700 28.800 ;
        RECT 78.200 28.200 78.500 28.800 ;
        RECT 80.600 28.200 80.900 33.800 ;
        RECT 81.400 29.800 81.800 30.200 ;
        RECT 78.200 27.800 78.600 28.200 ;
        RECT 79.000 27.800 79.400 28.200 ;
        RECT 80.600 27.800 81.000 28.200 ;
        RECT 79.000 27.100 79.300 27.800 ;
        RECT 77.400 26.800 79.300 27.100 ;
        RECT 81.400 27.200 81.700 29.800 ;
        RECT 82.200 29.200 82.500 33.800 ;
        RECT 82.200 28.800 82.600 29.200 ;
        RECT 83.000 28.200 83.300 33.800 ;
        RECT 87.000 33.200 87.300 35.800 ;
        RECT 90.200 35.200 90.500 35.800 ;
        RECT 91.800 35.200 92.100 38.800 ;
        RECT 94.200 37.800 94.600 38.200 ;
        RECT 92.600 35.800 93.000 36.200 ;
        RECT 92.600 35.200 92.900 35.800 ;
        RECT 88.600 34.800 89.000 35.200 ;
        RECT 90.200 34.800 90.600 35.200 ;
        RECT 91.000 34.800 91.400 35.200 ;
        RECT 91.800 34.800 92.200 35.200 ;
        RECT 92.600 34.800 93.000 35.200 ;
        RECT 88.600 34.200 88.900 34.800 ;
        RECT 91.000 34.200 91.300 34.800 ;
        RECT 88.600 33.800 89.000 34.200 ;
        RECT 91.000 33.800 91.400 34.200 ;
        RECT 91.800 33.800 92.200 34.200 ;
        RECT 83.800 33.100 84.200 33.200 ;
        RECT 84.600 33.100 85.000 33.200 ;
        RECT 83.800 32.800 85.000 33.100 ;
        RECT 87.000 32.800 87.400 33.200 ;
        RECT 88.600 33.100 89.000 33.200 ;
        RECT 89.400 33.100 89.800 33.200 ;
        RECT 88.600 32.800 89.800 33.100 ;
        RECT 87.000 30.200 87.300 32.800 ;
        RECT 87.800 31.800 88.200 32.200 ;
        RECT 87.000 29.800 87.400 30.200 ;
        RECT 86.200 28.800 86.600 29.200 ;
        RECT 86.200 28.200 86.500 28.800 ;
        RECT 83.000 27.800 83.400 28.200 ;
        RECT 83.800 27.800 84.200 28.200 ;
        RECT 86.200 27.800 86.600 28.200 ;
        RECT 83.800 27.200 84.100 27.800 ;
        RECT 87.800 27.200 88.100 31.800 ;
        RECT 91.800 28.200 92.100 33.800 ;
        RECT 94.200 33.200 94.500 37.800 ;
        RECT 95.800 36.800 96.200 37.200 ;
        RECT 95.800 35.200 96.100 36.800 ;
        RECT 95.800 34.800 96.200 35.200 ;
        RECT 96.600 34.100 96.900 42.800 ;
        RECT 97.400 36.200 97.700 45.800 ;
        RECT 99.000 45.200 99.300 45.800 ;
        RECT 99.800 45.200 100.100 45.800 ;
        RECT 101.400 45.200 101.700 45.800 ;
        RECT 105.400 45.200 105.700 48.800 ;
        RECT 107.800 47.800 108.200 48.200 ;
        RECT 107.800 47.200 108.100 47.800 ;
        RECT 108.600 47.200 108.900 51.800 ;
        RECT 106.200 47.100 106.600 47.200 ;
        RECT 107.000 47.100 107.400 47.200 ;
        RECT 106.200 46.800 107.400 47.100 ;
        RECT 107.800 46.800 108.200 47.200 ;
        RECT 108.600 46.800 109.000 47.200 ;
        RECT 106.200 45.800 106.600 46.200 ;
        RECT 108.600 45.800 109.000 46.200 ;
        RECT 99.000 44.800 99.400 45.200 ;
        RECT 99.800 44.800 100.200 45.200 ;
        RECT 101.400 44.800 101.800 45.200 ;
        RECT 104.600 44.800 105.000 45.200 ;
        RECT 105.400 44.800 105.800 45.200 ;
        RECT 104.600 43.200 104.900 44.800 ;
        RECT 106.200 44.200 106.500 45.800 ;
        RECT 108.600 45.200 108.900 45.800 ;
        RECT 108.600 44.800 109.000 45.200 ;
        RECT 106.200 43.800 106.600 44.200 ;
        RECT 104.600 42.800 105.000 43.200 ;
        RECT 102.200 41.800 102.600 42.200 ;
        RECT 108.600 41.800 109.000 42.200 ;
        RECT 101.400 36.800 101.800 37.200 ;
        RECT 97.400 35.800 97.800 36.200 ;
        RECT 101.400 35.200 101.700 36.800 ;
        RECT 101.400 34.800 101.800 35.200 ;
        RECT 95.800 33.800 96.900 34.100 ;
        RECT 102.200 34.200 102.500 41.800 ;
        RECT 108.600 40.200 108.900 41.800 ;
        RECT 108.600 39.800 109.000 40.200 ;
        RECT 104.600 38.100 105.000 38.200 ;
        RECT 105.400 38.100 105.800 38.200 ;
        RECT 104.600 37.800 105.800 38.100 ;
        RECT 107.800 38.100 108.200 38.200 ;
        RECT 108.600 38.100 109.000 38.200 ;
        RECT 107.800 37.800 109.000 38.100 ;
        RECT 104.600 36.800 105.000 37.200 ;
        RECT 106.200 36.800 106.600 37.200 ;
        RECT 104.600 36.200 104.900 36.800 ;
        RECT 103.000 35.800 103.400 36.200 ;
        RECT 104.600 35.800 105.000 36.200 ;
        RECT 103.000 35.200 103.300 35.800 ;
        RECT 103.000 34.800 103.400 35.200 ;
        RECT 104.600 34.800 105.000 35.200 ;
        RECT 104.600 34.200 104.900 34.800 ;
        RECT 106.200 34.200 106.500 36.800 ;
        RECT 107.000 36.100 107.400 36.200 ;
        RECT 107.800 36.100 108.200 36.200 ;
        RECT 107.000 35.800 108.200 36.100 ;
        RECT 108.600 35.800 109.000 36.200 ;
        RECT 102.200 33.800 102.600 34.200 ;
        RECT 104.600 33.800 105.000 34.200 ;
        RECT 106.200 33.800 106.600 34.200 ;
        RECT 108.600 34.100 108.900 35.800 ;
        RECT 109.400 35.200 109.700 52.800 ;
        RECT 115.000 51.800 115.400 52.200 ;
        RECT 113.400 50.800 113.800 51.200 ;
        RECT 113.400 49.200 113.700 50.800 ;
        RECT 111.800 48.800 112.200 49.200 ;
        RECT 113.400 48.800 113.800 49.200 ;
        RECT 111.800 48.200 112.100 48.800 ;
        RECT 111.800 47.800 112.200 48.200 ;
        RECT 112.600 47.800 113.000 48.200 ;
        RECT 110.200 46.800 110.600 47.200 ;
        RECT 110.200 45.200 110.500 46.800 ;
        RECT 110.200 44.800 110.600 45.200 ;
        RECT 111.000 41.800 111.400 42.200 ;
        RECT 110.200 37.800 110.600 38.200 ;
        RECT 110.200 35.200 110.500 37.800 ;
        RECT 111.000 36.200 111.300 41.800 ;
        RECT 112.600 39.200 112.900 47.800 ;
        RECT 115.000 47.200 115.300 51.800 ;
        RECT 115.000 46.800 115.400 47.200 ;
        RECT 115.000 46.200 115.300 46.800 ;
        RECT 115.800 46.200 116.100 53.800 ;
        RECT 119.000 53.200 119.300 53.800 ;
        RECT 119.000 52.800 119.400 53.200 ;
        RECT 123.000 52.800 123.400 53.200 ;
        RECT 125.400 52.800 125.800 53.200 ;
        RECT 126.200 52.800 126.600 53.200 ;
        RECT 117.400 47.100 117.800 47.200 ;
        RECT 118.200 47.100 118.600 47.200 ;
        RECT 117.400 46.800 118.600 47.100 ;
        RECT 119.000 46.200 119.300 52.800 ;
        RECT 119.800 51.800 120.200 52.200 ;
        RECT 115.000 45.800 115.400 46.200 ;
        RECT 115.800 45.800 116.200 46.200 ;
        RECT 119.000 45.800 119.400 46.200 ;
        RECT 115.800 45.200 116.100 45.800 ;
        RECT 115.800 44.800 116.200 45.200 ;
        RECT 117.400 44.800 117.800 45.200 ;
        RECT 119.800 45.100 120.100 51.800 ;
        RECT 123.000 49.200 123.300 52.800 ;
        RECT 125.400 52.200 125.700 52.800 ;
        RECT 125.400 51.800 125.800 52.200 ;
        RECT 126.200 51.100 126.500 52.800 ;
        RECT 125.400 50.800 126.500 51.100 ;
        RECT 129.400 51.800 129.800 52.200 ;
        RECT 123.000 48.800 123.400 49.200 ;
        RECT 120.600 47.100 121.000 47.200 ;
        RECT 121.400 47.100 121.800 47.200 ;
        RECT 120.600 46.800 121.800 47.100 ;
        RECT 123.000 46.800 123.400 47.200 ;
        RECT 124.600 46.800 125.000 47.200 ;
        RECT 125.400 47.100 125.700 50.800 ;
        RECT 126.200 48.800 126.600 49.200 ;
        RECT 127.000 48.800 127.400 49.200 ;
        RECT 126.200 48.200 126.500 48.800 ;
        RECT 126.200 47.800 126.600 48.200 ;
        RECT 126.200 47.100 126.600 47.200 ;
        RECT 125.400 46.800 126.600 47.100 ;
        RECT 121.400 46.100 121.800 46.200 ;
        RECT 122.200 46.100 122.600 46.200 ;
        RECT 121.400 45.800 122.600 46.100 ;
        RECT 123.000 45.200 123.300 46.800 ;
        RECT 124.600 46.200 124.900 46.800 ;
        RECT 127.000 46.200 127.300 48.800 ;
        RECT 129.400 47.200 129.700 51.800 ;
        RECT 131.800 47.200 132.100 53.800 ;
        RECT 136.600 52.100 137.000 52.200 ;
        RECT 137.400 52.100 137.800 52.200 ;
        RECT 136.600 51.800 137.800 52.100 ;
        RECT 138.200 49.800 138.600 50.200 ;
        RECT 138.200 49.200 138.500 49.800 ;
        RECT 138.200 48.800 138.600 49.200 ;
        RECT 134.200 48.100 134.600 48.200 ;
        RECT 135.000 48.100 135.400 48.200 ;
        RECT 139.000 48.100 139.300 54.800 ;
        RECT 134.200 47.800 135.400 48.100 ;
        RECT 138.200 47.800 139.300 48.100 ;
        RECT 139.800 48.200 140.100 65.800 ;
        RECT 140.600 64.800 141.000 65.200 ;
        RECT 140.600 64.200 140.900 64.800 ;
        RECT 140.600 63.800 141.000 64.200 ;
        RECT 141.400 54.200 141.700 65.800 ;
        RECT 142.200 63.800 142.600 64.200 ;
        RECT 142.200 63.200 142.500 63.800 ;
        RECT 142.200 62.800 142.600 63.200 ;
        RECT 145.400 62.200 145.700 66.800 ;
        RECT 147.000 64.200 147.300 67.800 ;
        RECT 148.600 67.200 148.900 71.800 ;
        RECT 148.600 66.800 149.000 67.200 ;
        RECT 149.400 66.200 149.700 81.800 ;
        RECT 150.200 76.200 150.500 82.800 ;
        RECT 150.200 75.800 150.600 76.200 ;
        RECT 149.400 65.800 149.800 66.200 ;
        RECT 147.000 63.800 147.400 64.200 ;
        RECT 145.400 61.800 145.800 62.200 ;
        RECT 143.800 59.100 144.200 59.200 ;
        RECT 144.600 59.100 145.000 59.200 ;
        RECT 143.800 58.800 145.000 59.100 ;
        RECT 144.600 55.100 145.000 55.200 ;
        RECT 145.400 55.100 145.800 55.200 ;
        RECT 144.600 54.800 145.800 55.100 ;
        RECT 146.200 55.100 146.600 55.200 ;
        RECT 147.000 55.100 147.400 55.200 ;
        RECT 146.200 54.800 147.400 55.100 ;
        RECT 149.400 55.100 149.800 55.200 ;
        RECT 150.200 55.100 150.600 55.200 ;
        RECT 149.400 54.800 150.600 55.100 ;
        RECT 141.400 53.800 141.800 54.200 ;
        RECT 142.200 54.100 142.600 54.200 ;
        RECT 143.000 54.100 143.400 54.200 ;
        RECT 142.200 53.800 143.400 54.100 ;
        RECT 148.600 53.800 149.000 54.200 ;
        RECT 148.600 53.200 148.900 53.800 ;
        RECT 142.200 52.800 142.600 53.200 ;
        RECT 143.000 52.800 143.400 53.200 ;
        RECT 147.800 52.800 148.200 53.200 ;
        RECT 148.600 52.800 149.000 53.200 ;
        RECT 142.200 52.200 142.500 52.800 ;
        RECT 142.200 51.800 142.600 52.200 ;
        RECT 141.400 50.800 141.800 51.200 ;
        RECT 141.400 49.200 141.700 50.800 ;
        RECT 141.400 48.800 141.800 49.200 ;
        RECT 139.800 47.800 140.200 48.200 ;
        RECT 129.400 46.800 129.800 47.200 ;
        RECT 131.800 46.800 132.200 47.200 ;
        RECT 134.200 47.100 134.600 47.200 ;
        RECT 135.000 47.100 135.400 47.200 ;
        RECT 134.200 46.800 135.400 47.100 ;
        RECT 136.600 46.800 137.000 47.200 ;
        RECT 123.800 45.800 124.200 46.200 ;
        RECT 124.600 45.800 125.000 46.200 ;
        RECT 127.000 45.800 127.400 46.200 ;
        RECT 127.800 46.100 128.200 46.200 ;
        RECT 128.600 46.100 129.000 46.200 ;
        RECT 127.800 45.800 129.000 46.100 ;
        RECT 120.600 45.100 121.000 45.200 ;
        RECT 119.800 44.800 121.000 45.100 ;
        RECT 121.400 44.800 121.800 45.200 ;
        RECT 123.000 44.800 123.400 45.200 ;
        RECT 117.400 43.200 117.700 44.800 ;
        RECT 117.400 42.800 117.800 43.200 ;
        RECT 115.800 41.800 116.200 42.200 ;
        RECT 113.400 39.800 113.800 40.200 ;
        RECT 112.600 38.800 113.000 39.200 ;
        RECT 111.000 35.800 111.400 36.200 ;
        RECT 113.400 35.200 113.700 39.800 ;
        RECT 115.800 35.200 116.100 41.800 ;
        RECT 117.400 37.200 117.700 42.800 ;
        RECT 121.400 40.200 121.700 44.800 ;
        RECT 123.000 44.200 123.300 44.800 ;
        RECT 123.000 43.800 123.400 44.200 ;
        RECT 123.800 41.200 124.100 45.800 ;
        RECT 123.800 40.800 124.200 41.200 ;
        RECT 127.000 40.800 127.400 41.200 ;
        RECT 121.400 39.800 121.800 40.200 ;
        RECT 117.400 36.800 117.800 37.200 ;
        RECT 118.200 36.100 118.600 36.200 ;
        RECT 117.400 35.800 118.600 36.100 ;
        RECT 120.600 35.800 121.000 36.200 ;
        RECT 109.400 34.800 109.800 35.200 ;
        RECT 110.200 34.800 110.600 35.200 ;
        RECT 111.800 34.800 112.200 35.200 ;
        RECT 113.400 34.800 113.800 35.200 ;
        RECT 115.000 34.800 115.400 35.200 ;
        RECT 115.800 34.800 116.200 35.200 ;
        RECT 111.800 34.200 112.100 34.800 ;
        RECT 109.400 34.100 109.800 34.200 ;
        RECT 108.600 33.800 109.800 34.100 ;
        RECT 111.800 33.800 112.200 34.200 ;
        RECT 112.600 33.800 113.000 34.200 ;
        RECT 115.000 34.100 115.300 34.800 ;
        RECT 115.800 34.100 116.200 34.200 ;
        RECT 115.000 33.800 116.200 34.100 ;
        RECT 94.200 32.800 94.600 33.200 ;
        RECT 95.800 29.200 96.100 33.800 ;
        RECT 98.200 32.800 98.600 33.200 ;
        RECT 111.000 33.100 111.400 33.200 ;
        RECT 111.800 33.100 112.200 33.200 ;
        RECT 111.000 32.800 112.200 33.100 ;
        RECT 98.200 32.200 98.500 32.800 ;
        RECT 97.400 31.800 97.800 32.200 ;
        RECT 98.200 31.800 98.600 32.200 ;
        RECT 99.000 31.800 99.400 32.200 ;
        RECT 111.000 31.800 111.400 32.200 ;
        RECT 95.800 28.800 96.200 29.200 ;
        RECT 97.400 28.200 97.700 31.800 ;
        RECT 99.000 30.200 99.300 31.800 ;
        RECT 99.000 29.800 99.400 30.200 ;
        RECT 103.800 29.800 104.200 30.200 ;
        RECT 103.800 29.200 104.100 29.800 ;
        RECT 111.000 29.200 111.300 31.800 ;
        RECT 112.600 30.200 112.900 33.800 ;
        RECT 115.000 31.800 115.400 32.200 ;
        RECT 112.600 29.800 113.000 30.200 ;
        RECT 115.000 29.200 115.300 31.800 ;
        RECT 117.400 29.200 117.700 35.800 ;
        RECT 119.000 35.100 119.400 35.200 ;
        RECT 119.800 35.100 120.200 35.200 ;
        RECT 119.000 34.800 120.200 35.100 ;
        RECT 119.000 33.800 119.400 34.200 ;
        RECT 118.200 32.800 118.600 33.200 ;
        RECT 118.200 32.200 118.500 32.800 ;
        RECT 118.200 31.800 118.600 32.200 ;
        RECT 119.000 30.200 119.300 33.800 ;
        RECT 120.600 31.200 120.900 35.800 ;
        RECT 123.800 35.100 124.200 35.200 ;
        RECT 124.600 35.100 125.000 35.200 ;
        RECT 123.800 34.800 125.000 35.100 ;
        RECT 122.200 33.800 122.600 34.200 ;
        RECT 121.400 32.800 121.800 33.200 ;
        RECT 121.400 31.200 121.700 32.800 ;
        RECT 120.600 30.800 121.000 31.200 ;
        RECT 121.400 30.800 121.800 31.200 ;
        RECT 122.200 30.200 122.500 33.800 ;
        RECT 127.000 33.200 127.300 40.800 ;
        RECT 128.600 38.800 129.000 39.200 ;
        RECT 128.600 38.200 128.900 38.800 ;
        RECT 128.600 37.800 129.000 38.200 ;
        RECT 129.400 33.200 129.700 46.800 ;
        RECT 130.200 45.800 130.600 46.200 ;
        RECT 131.000 45.800 131.400 46.200 ;
        RECT 130.200 45.200 130.500 45.800 ;
        RECT 130.200 44.800 130.600 45.200 ;
        RECT 131.000 43.200 131.300 45.800 ;
        RECT 131.800 45.200 132.100 46.800 ;
        RECT 136.600 46.200 136.900 46.800 ;
        RECT 136.600 45.800 137.000 46.200 ;
        RECT 131.800 44.800 132.200 45.200 ;
        RECT 136.600 44.800 137.000 45.200 ;
        RECT 136.600 44.200 136.900 44.800 ;
        RECT 136.600 43.800 137.000 44.200 ;
        RECT 131.000 42.800 131.400 43.200 ;
        RECT 138.200 42.200 138.500 47.800 ;
        RECT 139.800 47.200 140.100 47.800 ;
        RECT 139.800 46.800 140.200 47.200 ;
        RECT 140.600 46.800 141.000 47.200 ;
        RECT 139.800 45.800 140.200 46.200 ;
        RECT 139.800 45.200 140.100 45.800 ;
        RECT 139.800 44.800 140.200 45.200 ;
        RECT 131.000 41.800 131.400 42.200 ;
        RECT 133.400 41.800 133.800 42.200 ;
        RECT 138.200 41.800 138.600 42.200 ;
        RECT 127.000 32.800 127.400 33.200 ;
        RECT 129.400 32.800 129.800 33.200 ;
        RECT 119.000 29.800 119.400 30.200 ;
        RECT 122.200 29.800 122.600 30.200 ;
        RECT 103.800 28.800 104.200 29.200 ;
        RECT 111.000 28.800 111.400 29.200 ;
        RECT 114.200 28.800 114.600 29.200 ;
        RECT 115.000 28.800 115.400 29.200 ;
        RECT 117.400 28.800 117.800 29.200 ;
        RECT 121.400 28.800 121.800 29.200 ;
        RECT 114.200 28.200 114.500 28.800 ;
        RECT 91.800 27.800 92.200 28.200 ;
        RECT 93.400 27.800 93.800 28.200 ;
        RECT 95.800 28.100 96.200 28.200 ;
        RECT 96.600 28.100 97.000 28.200 ;
        RECT 95.800 27.800 97.000 28.100 ;
        RECT 97.400 27.800 97.800 28.200 ;
        RECT 105.400 27.800 105.800 28.200 ;
        RECT 110.200 27.800 110.600 28.200 ;
        RECT 111.800 27.800 112.200 28.200 ;
        RECT 114.200 27.800 114.600 28.200 ;
        RECT 115.000 28.100 115.400 28.200 ;
        RECT 115.800 28.100 116.200 28.200 ;
        RECT 118.200 28.100 118.600 28.200 ;
        RECT 115.000 27.800 116.200 28.100 ;
        RECT 117.400 27.800 118.600 28.100 ;
        RECT 81.400 26.800 81.800 27.200 ;
        RECT 83.800 26.800 84.200 27.200 ;
        RECT 87.800 26.800 88.200 27.200 ;
        RECT 89.400 26.800 89.800 27.200 ;
        RECT 75.800 26.200 76.100 26.800 ;
        RECT 89.400 26.200 89.700 26.800 ;
        RECT 91.800 26.200 92.100 27.800 ;
        RECT 92.600 26.800 93.000 27.200 ;
        RECT 92.600 26.200 92.900 26.800 ;
        RECT 71.000 25.800 71.400 26.200 ;
        RECT 75.000 25.800 75.400 26.200 ;
        RECT 75.800 25.800 76.200 26.200 ;
        RECT 76.600 25.800 77.000 26.200 ;
        RECT 80.600 25.800 81.000 26.200 ;
        RECT 89.400 25.800 89.800 26.200 ;
        RECT 91.800 25.800 92.200 26.200 ;
        RECT 92.600 25.800 93.000 26.200 ;
        RECT 93.400 26.100 93.700 27.800 ;
        RECT 105.400 27.200 105.700 27.800 ;
        RECT 110.200 27.200 110.500 27.800 ;
        RECT 111.800 27.200 112.100 27.800 ;
        RECT 94.200 27.100 94.600 27.200 ;
        RECT 95.000 27.100 95.400 27.200 ;
        RECT 94.200 26.800 95.400 27.100 ;
        RECT 97.400 27.100 97.800 27.200 ;
        RECT 98.200 27.100 98.600 27.200 ;
        RECT 97.400 26.800 98.600 27.100 ;
        RECT 99.800 27.100 100.200 27.200 ;
        RECT 100.600 27.100 101.000 27.200 ;
        RECT 99.800 26.800 101.000 27.100 ;
        RECT 101.400 26.800 101.800 27.200 ;
        RECT 102.200 26.900 102.600 27.000 ;
        RECT 103.000 26.900 103.400 27.000 ;
        RECT 94.200 26.100 94.600 26.200 ;
        RECT 93.400 25.800 94.600 26.100 ;
        RECT 99.000 25.800 99.400 26.200 ;
        RECT 71.000 25.200 71.300 25.800 ;
        RECT 76.600 25.200 76.900 25.800 ;
        RECT 71.000 24.800 71.400 25.200 ;
        RECT 75.800 24.800 76.200 25.200 ;
        RECT 76.600 24.800 77.000 25.200 ;
        RECT 74.200 18.800 74.600 19.200 ;
        RECT 74.200 18.200 74.500 18.800 ;
        RECT 72.600 17.800 73.000 18.200 ;
        RECT 74.200 17.800 74.600 18.200 ;
        RECT 72.600 16.200 72.900 17.800 ;
        RECT 74.200 17.100 74.600 17.200 ;
        RECT 75.000 17.100 75.400 17.200 ;
        RECT 74.200 16.800 75.400 17.100 ;
        RECT 72.600 15.800 73.000 16.200 ;
        RECT 75.000 15.800 75.400 16.200 ;
        RECT 75.000 15.200 75.300 15.800 ;
        RECT 66.200 15.100 66.600 15.200 ;
        RECT 67.000 15.100 67.400 15.200 ;
        RECT 66.200 14.800 67.400 15.100 ;
        RECT 67.800 14.800 68.200 15.200 ;
        RECT 70.200 14.800 70.600 15.200 ;
        RECT 72.600 14.800 73.000 15.200 ;
        RECT 75.000 14.800 75.400 15.200 ;
        RECT 70.200 14.200 70.500 14.800 ;
        RECT 72.600 14.200 72.900 14.800 ;
        RECT 70.200 13.800 70.600 14.200 ;
        RECT 72.600 13.800 73.000 14.200 ;
        RECT 65.400 12.800 65.800 13.200 ;
        RECT 68.600 12.100 69.000 12.200 ;
        RECT 69.400 12.100 69.800 12.200 ;
        RECT 68.600 11.800 69.800 12.100 ;
        RECT 64.600 10.800 65.000 11.200 ;
        RECT 64.600 9.200 64.900 10.800 ;
        RECT 66.200 9.800 66.600 10.200 ;
        RECT 66.200 9.200 66.500 9.800 ;
        RECT 58.200 8.800 58.600 9.200 ;
        RECT 61.400 8.800 61.800 9.200 ;
        RECT 63.800 8.800 64.200 9.200 ;
        RECT 64.600 8.800 65.000 9.200 ;
        RECT 66.200 8.800 66.600 9.200 ;
        RECT 71.000 9.100 71.400 9.200 ;
        RECT 71.800 9.100 72.200 9.200 ;
        RECT 71.000 8.800 72.200 9.100 ;
        RECT 75.800 8.200 76.100 24.800 ;
        RECT 80.600 23.200 80.900 25.800 ;
        RECT 85.400 25.100 85.800 25.200 ;
        RECT 86.200 25.100 86.600 25.200 ;
        RECT 85.400 24.800 86.600 25.100 ;
        RECT 87.000 24.800 87.400 25.200 ;
        RECT 80.600 22.800 81.000 23.200 ;
        RECT 80.600 22.200 80.900 22.800 ;
        RECT 77.400 21.800 77.800 22.200 ;
        RECT 80.600 21.800 81.000 22.200 ;
        RECT 77.400 20.200 77.700 21.800 ;
        RECT 79.800 20.800 80.200 21.200 ;
        RECT 77.400 19.800 77.800 20.200 ;
        RECT 79.800 19.200 80.100 20.800 ;
        RECT 79.800 18.800 80.200 19.200 ;
        RECT 76.600 16.100 77.000 16.200 ;
        RECT 77.400 16.100 77.800 16.200 ;
        RECT 76.600 15.800 77.800 16.100 ;
        RECT 81.300 15.900 81.700 16.300 ;
        RECT 84.600 15.900 85.000 16.300 ;
        RECT 76.600 13.800 77.000 14.200 ;
        RECT 76.600 13.200 76.900 13.800 ;
        RECT 81.300 13.500 81.600 15.900 ;
        RECT 82.600 14.200 83.000 14.300 ;
        RECT 84.700 14.200 85.000 15.900 ;
        RECT 85.400 16.100 85.800 16.200 ;
        RECT 86.200 16.100 86.600 16.200 ;
        RECT 85.400 15.800 86.600 16.100 ;
        RECT 86.200 14.800 86.600 15.200 ;
        RECT 82.600 13.900 85.000 14.200 ;
        RECT 82.200 13.500 82.600 13.600 ;
        RECT 83.900 13.500 84.300 13.600 ;
        RECT 84.700 13.500 85.000 13.900 ;
        RECT 76.600 12.800 77.000 13.200 ;
        RECT 81.300 13.100 81.700 13.500 ;
        RECT 82.200 13.200 84.300 13.500 ;
        RECT 82.200 9.200 82.500 13.200 ;
        RECT 84.600 13.100 85.000 13.500 ;
        RECT 85.400 13.800 85.800 14.200 ;
        RECT 85.400 11.200 85.700 13.800 ;
        RECT 86.200 13.200 86.500 14.800 ;
        RECT 86.200 12.800 86.600 13.200 ;
        RECT 86.200 11.800 86.600 12.200 ;
        RECT 83.000 10.800 83.400 11.200 ;
        RECT 85.400 10.800 85.800 11.200 ;
        RECT 83.000 9.200 83.300 10.800 ;
        RECT 86.200 9.200 86.500 11.800 ;
        RECT 87.000 9.200 87.300 24.800 ;
        RECT 92.600 24.100 93.000 24.200 ;
        RECT 92.600 23.800 93.700 24.100 ;
        RECT 88.600 21.800 89.000 22.200 ;
        RECT 87.800 15.800 88.200 16.200 ;
        RECT 87.800 15.200 88.100 15.800 ;
        RECT 87.800 14.800 88.200 15.200 ;
        RECT 88.600 14.200 88.900 21.800 ;
        RECT 93.400 19.200 93.700 23.800 ;
        RECT 94.200 23.200 94.500 25.800 ;
        RECT 99.000 25.200 99.300 25.800 ;
        RECT 99.000 24.800 99.400 25.200 ;
        RECT 94.200 22.800 94.600 23.200 ;
        RECT 93.400 18.800 93.800 19.200 ;
        RECT 94.200 17.800 94.600 18.200 ;
        RECT 98.200 17.800 98.600 18.200 ;
        RECT 94.200 16.200 94.500 17.800 ;
        RECT 95.800 16.800 96.200 17.200 ;
        RECT 94.200 15.800 94.600 16.200 ;
        RECT 95.800 15.200 96.100 16.800 ;
        RECT 90.200 14.800 90.600 15.200 ;
        RECT 91.000 14.800 91.400 15.200 ;
        RECT 95.800 14.800 96.200 15.200 ;
        RECT 90.200 14.200 90.500 14.800 ;
        RECT 91.000 14.200 91.300 14.800 ;
        RECT 88.600 13.800 89.000 14.200 ;
        RECT 89.400 13.800 89.800 14.200 ;
        RECT 90.200 13.800 90.600 14.200 ;
        RECT 91.000 13.800 91.400 14.200 ;
        RECT 91.800 13.800 92.200 14.200 ;
        RECT 89.400 11.200 89.700 13.800 ;
        RECT 91.800 13.200 92.100 13.800 ;
        RECT 91.800 12.800 92.200 13.200 ;
        RECT 94.200 12.800 94.600 13.200 ;
        RECT 89.400 10.800 89.800 11.200 ;
        RECT 78.200 8.800 78.600 9.200 ;
        RECT 81.400 8.800 81.800 9.200 ;
        RECT 82.200 8.800 82.600 9.200 ;
        RECT 83.000 8.800 83.400 9.200 ;
        RECT 86.200 8.800 86.600 9.200 ;
        RECT 87.000 8.800 87.400 9.200 ;
        RECT 78.200 8.200 78.500 8.800 ;
        RECT 69.400 8.100 69.800 8.200 ;
        RECT 70.200 8.100 70.600 8.200 ;
        RECT 69.400 7.800 70.600 8.100 ;
        RECT 75.800 7.800 76.200 8.200 ;
        RECT 78.200 7.800 78.600 8.200 ;
        RECT 75.800 7.200 76.100 7.800 ;
        RECT 53.400 7.100 53.800 7.200 ;
        RECT 54.200 7.100 54.600 7.200 ;
        RECT 53.400 6.800 54.600 7.100 ;
        RECT 55.800 7.100 56.200 7.200 ;
        RECT 56.600 7.100 57.000 7.200 ;
        RECT 55.800 6.800 57.000 7.100 ;
        RECT 75.800 6.800 76.200 7.200 ;
        RECT 79.000 7.100 79.400 7.200 ;
        RECT 79.800 7.100 80.200 7.200 ;
        RECT 79.000 6.800 80.200 7.100 ;
        RECT 36.600 6.100 37.000 6.200 ;
        RECT 37.400 6.100 37.800 6.200 ;
        RECT 36.600 5.800 37.800 6.100 ;
        RECT 39.800 5.800 40.200 6.200 ;
        RECT 47.800 6.100 48.200 6.200 ;
        RECT 48.600 6.100 49.000 6.200 ;
        RECT 47.800 5.800 49.000 6.100 ;
        RECT 49.400 5.800 49.800 6.200 ;
        RECT 52.600 5.800 53.000 6.200 ;
        RECT 70.200 6.100 70.600 6.200 ;
        RECT 71.000 6.100 71.400 6.200 ;
        RECT 70.200 5.800 71.400 6.100 ;
        RECT 73.400 6.100 73.800 6.200 ;
        RECT 74.200 6.100 74.600 6.200 ;
        RECT 73.400 5.800 74.600 6.100 ;
        RECT 79.000 6.100 79.400 6.200 ;
        RECT 79.800 6.100 80.200 6.200 ;
        RECT 79.000 5.800 80.200 6.100 ;
        RECT 29.500 4.700 29.900 5.100 ;
        RECT 30.200 4.800 31.400 5.100 ;
        RECT 32.600 4.700 33.000 5.100 ;
        RECT 39.800 5.200 40.100 5.800 ;
        RECT 81.400 5.200 81.700 8.800 ;
        RECT 82.200 7.800 82.600 8.200 ;
        RECT 84.600 7.800 85.000 8.200 ;
        RECT 86.200 7.800 86.600 8.200 ;
        RECT 91.000 7.800 91.400 8.200 ;
        RECT 82.200 6.200 82.500 7.800 ;
        RECT 84.600 7.200 84.900 7.800 ;
        RECT 86.200 7.200 86.500 7.800 ;
        RECT 91.000 7.200 91.300 7.800 ;
        RECT 94.200 7.200 94.500 12.800 ;
        RECT 95.800 9.100 96.200 9.200 ;
        RECT 96.600 9.100 97.000 9.200 ;
        RECT 95.800 8.800 97.000 9.100 ;
        RECT 98.200 7.200 98.500 17.800 ;
        RECT 101.400 15.200 101.700 26.800 ;
        RECT 102.200 26.600 103.400 26.900 ;
        RECT 105.400 26.800 105.800 27.200 ;
        RECT 107.800 26.800 108.200 27.200 ;
        RECT 108.600 26.800 109.000 27.200 ;
        RECT 110.200 26.800 110.600 27.200 ;
        RECT 111.800 26.800 112.200 27.200 ;
        RECT 113.400 26.800 113.800 27.200 ;
        RECT 115.800 26.800 116.200 27.200 ;
        RECT 116.600 26.800 117.000 27.200 ;
        RECT 105.400 25.200 105.700 26.800 ;
        RECT 107.800 26.200 108.100 26.800 ;
        RECT 107.800 25.800 108.200 26.200 ;
        RECT 105.400 24.800 105.800 25.200 ;
        RECT 107.000 25.100 107.400 25.200 ;
        RECT 107.800 25.100 108.200 25.200 ;
        RECT 107.000 24.800 108.200 25.100 ;
        RECT 104.600 23.800 105.000 24.200 ;
        RECT 104.600 22.200 104.900 23.800 ;
        RECT 107.000 22.800 107.400 23.200 ;
        RECT 103.800 22.100 104.200 22.200 ;
        RECT 104.600 22.100 105.000 22.200 ;
        RECT 103.800 21.800 105.000 22.100 ;
        RECT 103.800 19.800 104.200 20.200 ;
        RECT 99.000 14.800 99.400 15.200 ;
        RECT 101.400 14.800 101.800 15.200 ;
        RECT 99.000 14.200 99.300 14.800 ;
        RECT 99.000 13.800 99.400 14.200 ;
        RECT 99.800 13.800 100.200 14.200 ;
        RECT 84.600 6.800 85.000 7.200 ;
        RECT 86.200 6.800 86.600 7.200 ;
        RECT 90.200 6.800 90.600 7.200 ;
        RECT 91.000 6.800 91.400 7.200 ;
        RECT 91.800 7.100 92.200 7.200 ;
        RECT 92.600 7.100 93.000 7.200 ;
        RECT 91.800 6.800 93.000 7.100 ;
        RECT 94.200 6.800 94.600 7.200 ;
        RECT 95.000 6.800 95.400 7.200 ;
        RECT 98.200 6.800 98.600 7.200 ;
        RECT 84.600 6.200 84.900 6.800 ;
        RECT 90.200 6.200 90.500 6.800 ;
        RECT 95.000 6.200 95.300 6.800 ;
        RECT 99.000 6.200 99.300 13.800 ;
        RECT 99.800 13.200 100.100 13.800 ;
        RECT 99.800 12.800 100.200 13.200 ;
        RECT 102.200 12.800 102.600 13.200 ;
        RECT 100.600 7.800 101.000 8.200 ;
        RECT 100.600 7.200 100.900 7.800 ;
        RECT 102.200 7.200 102.500 12.800 ;
        RECT 103.800 8.100 104.100 19.800 ;
        RECT 107.000 17.200 107.300 22.800 ;
        RECT 108.600 20.200 108.900 26.800 ;
        RECT 109.400 25.800 109.800 26.200 ;
        RECT 112.600 25.800 113.000 26.200 ;
        RECT 109.400 25.200 109.700 25.800 ;
        RECT 109.400 24.800 109.800 25.200 ;
        RECT 112.600 22.200 112.900 25.800 ;
        RECT 113.400 24.200 113.700 26.800 ;
        RECT 115.800 26.200 116.100 26.800 ;
        RECT 116.600 26.200 116.900 26.800 ;
        RECT 115.800 25.800 116.200 26.200 ;
        RECT 116.600 25.800 117.000 26.200 ;
        RECT 117.400 26.100 117.700 27.800 ;
        RECT 121.400 27.200 121.700 28.800 ;
        RECT 127.000 28.200 127.300 32.800 ;
        RECT 128.600 29.800 129.000 30.200 ;
        RECT 127.000 27.800 127.400 28.200 ;
        RECT 128.600 27.200 128.900 29.800 ;
        RECT 118.200 27.100 118.600 27.200 ;
        RECT 119.000 27.100 119.400 27.200 ;
        RECT 118.200 26.800 119.400 27.100 ;
        RECT 121.400 26.800 121.800 27.200 ;
        RECT 123.800 27.100 124.200 27.200 ;
        RECT 124.600 27.100 125.000 27.200 ;
        RECT 123.800 26.800 125.000 27.100 ;
        RECT 128.600 26.800 129.000 27.200 ;
        RECT 129.400 27.100 129.800 27.200 ;
        RECT 130.200 27.100 130.600 27.200 ;
        RECT 129.400 26.800 130.600 27.100 ;
        RECT 131.000 27.100 131.300 41.800 ;
        RECT 133.400 41.200 133.700 41.800 ;
        RECT 140.600 41.200 140.900 46.800 ;
        RECT 141.400 42.800 141.800 43.200 ;
        RECT 133.400 40.800 133.800 41.200 ;
        RECT 135.800 40.800 136.200 41.200 ;
        RECT 136.600 40.800 137.000 41.200 ;
        RECT 140.600 40.800 141.000 41.200 ;
        RECT 133.400 39.800 133.800 40.200 ;
        RECT 133.400 39.200 133.700 39.800 ;
        RECT 133.400 38.800 133.800 39.200 ;
        RECT 135.800 37.200 136.100 40.800 ;
        RECT 136.600 39.200 136.900 40.800 ;
        RECT 141.400 39.200 141.700 42.800 ;
        RECT 136.600 38.800 137.000 39.200 ;
        RECT 141.400 38.800 141.800 39.200 ;
        RECT 135.800 36.800 136.200 37.200 ;
        RECT 137.400 36.100 137.800 36.200 ;
        RECT 138.200 36.100 138.600 36.200 ;
        RECT 137.400 35.800 138.600 36.100 ;
        RECT 139.000 35.800 139.400 36.200 ;
        RECT 134.200 34.800 134.600 35.200 ;
        RECT 135.800 35.100 136.200 35.200 ;
        RECT 136.600 35.100 137.000 35.200 ;
        RECT 135.800 34.800 137.000 35.100 ;
        RECT 137.400 35.100 137.800 35.200 ;
        RECT 138.200 35.100 138.600 35.200 ;
        RECT 137.400 34.800 138.600 35.100 ;
        RECT 134.200 34.200 134.500 34.800 ;
        RECT 131.800 33.800 132.200 34.200 ;
        RECT 134.200 33.800 134.600 34.200 ;
        RECT 131.800 32.200 132.100 33.800 ;
        RECT 132.600 33.100 133.000 33.200 ;
        RECT 133.400 33.100 133.800 33.200 ;
        RECT 132.600 32.800 133.800 33.100 ;
        RECT 131.800 31.800 132.200 32.200 ;
        RECT 132.600 27.800 133.000 28.200 ;
        RECT 131.000 26.800 132.100 27.100 ;
        RECT 123.800 26.100 124.200 26.200 ;
        RECT 124.600 26.100 125.000 26.200 ;
        RECT 117.400 25.800 118.500 26.100 ;
        RECT 123.800 25.800 125.000 26.100 ;
        RECT 126.200 25.800 126.600 26.200 ;
        RECT 127.000 26.100 127.400 26.200 ;
        RECT 127.800 26.100 128.200 26.200 ;
        RECT 127.000 25.800 128.200 26.100 ;
        RECT 113.400 23.800 113.800 24.200 ;
        RECT 112.600 21.800 113.000 22.200 ;
        RECT 111.800 20.800 112.200 21.200 ;
        RECT 108.600 19.800 109.000 20.200 ;
        RECT 105.400 17.100 105.800 17.200 ;
        RECT 106.200 17.100 106.600 17.200 ;
        RECT 105.400 16.800 106.600 17.100 ;
        RECT 107.000 16.800 107.400 17.200 ;
        RECT 107.000 16.100 107.400 16.200 ;
        RECT 104.600 15.800 107.400 16.100 ;
        RECT 110.200 15.800 110.600 16.200 ;
        RECT 104.600 15.200 104.900 15.800 ;
        RECT 110.200 15.200 110.500 15.800 ;
        RECT 111.800 15.200 112.100 20.800 ;
        RECT 113.400 19.800 113.800 20.200 ;
        RECT 113.400 16.200 113.700 19.800 ;
        RECT 114.200 17.800 114.600 18.200 ;
        RECT 113.400 15.800 113.800 16.200 ;
        RECT 113.400 15.200 113.700 15.800 ;
        RECT 104.600 14.800 105.000 15.200 ;
        RECT 105.400 14.800 105.800 15.200 ;
        RECT 107.000 14.800 107.400 15.200 ;
        RECT 110.200 14.800 110.600 15.200 ;
        RECT 111.800 14.800 112.200 15.200 ;
        RECT 113.400 14.800 113.800 15.200 ;
        RECT 105.400 14.200 105.700 14.800 ;
        RECT 104.600 13.800 105.000 14.200 ;
        RECT 105.400 13.800 105.800 14.200 ;
        RECT 104.600 13.200 104.900 13.800 ;
        RECT 104.600 12.800 105.000 13.200 ;
        RECT 107.000 9.200 107.300 14.800 ;
        RECT 114.200 14.200 114.500 17.800 ;
        RECT 115.000 17.100 115.400 17.200 ;
        RECT 115.800 17.100 116.200 17.200 ;
        RECT 115.000 16.800 116.200 17.100 ;
        RECT 115.000 14.800 115.400 15.200 ;
        RECT 107.800 13.800 108.200 14.200 ;
        RECT 109.400 14.100 109.800 14.200 ;
        RECT 110.200 14.100 110.600 14.200 ;
        RECT 109.400 13.800 110.600 14.100 ;
        RECT 111.000 13.800 111.400 14.200 ;
        RECT 114.200 13.800 114.600 14.200 ;
        RECT 107.800 12.200 108.100 13.800 ;
        RECT 111.000 13.200 111.300 13.800 ;
        RECT 109.400 12.800 109.800 13.200 ;
        RECT 111.000 12.800 111.400 13.200 ;
        RECT 111.800 12.800 112.200 13.200 ;
        RECT 112.600 12.800 113.000 13.200 ;
        RECT 107.800 11.800 108.200 12.200 ;
        RECT 107.800 10.200 108.100 11.800 ;
        RECT 107.800 9.800 108.200 10.200 ;
        RECT 109.400 9.200 109.700 12.800 ;
        RECT 111.800 12.200 112.100 12.800 ;
        RECT 111.800 11.800 112.200 12.200 ;
        RECT 110.200 10.800 110.600 11.200 ;
        RECT 107.000 8.800 107.400 9.200 ;
        RECT 109.400 8.800 109.800 9.200 ;
        RECT 104.600 8.100 105.000 8.200 ;
        RECT 103.800 7.800 105.000 8.100 ;
        RECT 100.600 6.800 101.000 7.200 ;
        RECT 102.200 6.800 102.600 7.200 ;
        RECT 82.200 5.800 82.600 6.200 ;
        RECT 84.600 5.800 85.000 6.200 ;
        RECT 86.200 5.800 86.600 6.200 ;
        RECT 90.200 5.800 90.600 6.200 ;
        RECT 92.600 6.100 93.000 6.200 ;
        RECT 93.400 6.100 93.800 6.200 ;
        RECT 92.600 5.800 94.500 6.100 ;
        RECT 95.000 5.800 95.400 6.200 ;
        RECT 95.800 5.800 96.200 6.200 ;
        RECT 99.000 5.800 99.400 6.200 ;
        RECT 101.400 6.100 101.800 6.200 ;
        RECT 102.200 6.100 102.600 6.200 ;
        RECT 101.400 5.800 102.600 6.100 ;
        RECT 103.000 6.100 103.400 6.200 ;
        RECT 103.800 6.100 104.200 6.200 ;
        RECT 103.000 5.800 104.200 6.100 ;
        RECT 106.200 6.100 106.600 6.200 ;
        RECT 107.000 6.100 107.300 8.800 ;
        RECT 110.200 6.200 110.500 10.800 ;
        RECT 111.000 9.800 111.400 10.200 ;
        RECT 111.000 8.200 111.300 9.800 ;
        RECT 112.600 8.200 112.900 12.800 ;
        RECT 115.000 10.200 115.300 14.800 ;
        RECT 118.200 14.100 118.500 25.800 ;
        RECT 119.000 25.100 119.400 25.200 ;
        RECT 119.800 25.100 120.200 25.200 ;
        RECT 119.000 24.800 120.200 25.100 ;
        RECT 122.200 24.800 122.600 25.200 ;
        RECT 122.200 23.200 122.500 24.800 ;
        RECT 122.200 22.800 122.600 23.200 ;
        RECT 126.200 22.200 126.500 25.800 ;
        RECT 126.200 21.800 126.600 22.200 ;
        RECT 124.600 20.800 125.000 21.200 ;
        RECT 123.000 19.800 123.400 20.200 ;
        RECT 123.000 19.200 123.300 19.800 ;
        RECT 123.000 18.800 123.400 19.200 ;
        RECT 119.800 16.800 120.200 17.200 ;
        RECT 119.000 15.100 119.400 15.200 ;
        RECT 119.800 15.100 120.100 16.800 ;
        RECT 121.400 15.800 121.800 16.200 ;
        RECT 119.000 14.800 120.100 15.100 ;
        RECT 120.600 15.100 121.000 15.200 ;
        RECT 121.400 15.100 121.700 15.800 ;
        RECT 120.600 14.800 121.700 15.100 ;
        RECT 118.200 13.800 119.300 14.100 ;
        RECT 116.600 12.800 117.000 13.200 ;
        RECT 115.000 9.800 115.400 10.200 ;
        RECT 116.600 9.200 116.900 12.800 ;
        RECT 117.400 11.800 117.800 12.200 ;
        RECT 117.400 11.200 117.700 11.800 ;
        RECT 117.400 10.800 117.800 11.200 ;
        RECT 119.000 9.200 119.300 13.800 ;
        RECT 120.600 13.800 121.000 14.200 ;
        RECT 120.600 12.200 120.900 13.800 ;
        RECT 124.600 13.200 124.900 20.800 ;
        RECT 126.200 19.200 126.500 21.800 ;
        RECT 128.600 21.200 128.900 26.800 ;
        RECT 130.200 26.100 130.600 26.200 ;
        RECT 131.000 26.100 131.400 26.200 ;
        RECT 130.200 25.800 131.400 26.100 ;
        RECT 128.600 20.800 129.000 21.200 ;
        RECT 126.200 18.800 126.600 19.200 ;
        RECT 127.000 18.800 127.400 19.200 ;
        RECT 126.200 16.800 126.600 17.200 ;
        RECT 126.200 14.200 126.500 16.800 ;
        RECT 127.000 15.200 127.300 18.800 ;
        RECT 127.800 17.100 128.200 17.200 ;
        RECT 128.600 17.100 129.000 17.200 ;
        RECT 127.800 16.800 129.000 17.100 ;
        RECT 131.800 16.200 132.100 26.800 ;
        RECT 132.600 26.200 132.900 27.800 ;
        RECT 133.400 26.800 133.800 27.200 ;
        RECT 133.400 26.200 133.700 26.800 ;
        RECT 132.600 25.800 133.000 26.200 ;
        RECT 133.400 25.800 133.800 26.200 ;
        RECT 132.600 19.200 132.900 25.800 ;
        RECT 132.600 18.800 133.000 19.200 ;
        RECT 133.400 18.800 133.800 19.200 ;
        RECT 133.400 17.200 133.700 18.800 ;
        RECT 134.200 18.200 134.500 33.800 ;
        RECT 138.200 32.800 138.600 33.200 ;
        RECT 138.200 29.200 138.500 32.800 ;
        RECT 138.200 28.800 138.600 29.200 ;
        RECT 139.000 28.200 139.300 35.800 ;
        RECT 140.600 35.100 141.000 35.200 ;
        RECT 141.400 35.100 141.800 35.200 ;
        RECT 140.600 34.800 141.800 35.100 ;
        RECT 139.800 34.100 140.200 34.200 ;
        RECT 140.600 34.100 141.000 34.200 ;
        RECT 139.800 33.800 141.000 34.100 ;
        RECT 141.400 33.200 141.700 34.800 ;
        RECT 142.200 34.200 142.500 51.800 ;
        RECT 143.000 45.200 143.300 52.800 ;
        RECT 147.800 50.200 148.100 52.800 ;
        RECT 149.400 51.800 149.800 52.200 ;
        RECT 149.400 51.100 149.700 51.800 ;
        RECT 150.200 51.100 150.600 51.200 ;
        RECT 149.400 50.800 150.600 51.100 ;
        RECT 147.800 49.800 148.200 50.200 ;
        RECT 149.400 49.800 149.800 50.200 ;
        RECT 149.400 49.200 149.700 49.800 ;
        RECT 149.400 48.800 149.800 49.200 ;
        RECT 150.200 48.800 150.600 49.200 ;
        RECT 147.800 47.800 148.200 48.200 ;
        RECT 147.800 47.200 148.100 47.800 ;
        RECT 147.800 46.800 148.200 47.200 ;
        RECT 150.200 46.200 150.500 48.800 ;
        RECT 145.400 45.800 145.800 46.200 ;
        RECT 150.200 45.800 150.600 46.200 ;
        RECT 145.400 45.200 145.700 45.800 ;
        RECT 143.000 44.800 143.400 45.200 ;
        RECT 145.400 44.800 145.800 45.200 ;
        RECT 143.000 35.100 143.400 35.200 ;
        RECT 143.800 35.100 144.200 35.200 ;
        RECT 143.000 34.800 144.200 35.100 ;
        RECT 142.200 33.800 142.600 34.200 ;
        RECT 147.800 33.800 148.200 34.200 ;
        RECT 141.400 32.800 141.800 33.200 ;
        RECT 146.200 31.800 146.600 32.200 ;
        RECT 139.800 29.100 140.200 29.200 ;
        RECT 140.600 29.100 141.000 29.200 ;
        RECT 139.800 28.800 141.000 29.100 ;
        RECT 139.000 27.800 139.400 28.200 ;
        RECT 145.400 27.800 145.800 28.200 ;
        RECT 136.600 27.100 137.000 27.200 ;
        RECT 137.400 27.100 137.800 27.200 ;
        RECT 136.600 26.800 137.800 27.100 ;
        RECT 139.000 26.200 139.300 27.800 ;
        RECT 145.400 27.200 145.700 27.800 ;
        RECT 141.400 27.100 141.800 27.200 ;
        RECT 142.200 27.100 142.600 27.200 ;
        RECT 141.400 26.800 142.600 27.100 ;
        RECT 143.000 26.800 143.400 27.200 ;
        RECT 145.400 26.800 145.800 27.200 ;
        RECT 139.000 25.800 139.400 26.200 ;
        RECT 141.400 25.800 141.800 26.200 ;
        RECT 135.800 24.800 136.200 25.200 ;
        RECT 134.200 17.800 134.600 18.200 ;
        RECT 135.800 17.200 136.100 24.800 ;
        RECT 140.600 17.800 141.000 18.200 ;
        RECT 133.400 16.800 133.800 17.200 ;
        RECT 135.800 16.800 136.200 17.200 ;
        RECT 131.800 15.800 132.200 16.200 ;
        RECT 136.600 15.800 137.000 16.200 ;
        RECT 138.200 16.100 138.600 16.200 ;
        RECT 139.000 16.100 139.400 16.200 ;
        RECT 138.200 15.800 139.400 16.100 ;
        RECT 136.600 15.200 136.900 15.800 ;
        RECT 127.000 14.800 127.400 15.200 ;
        RECT 128.600 15.100 129.000 15.200 ;
        RECT 127.800 14.800 129.000 15.100 ;
        RECT 133.400 15.100 133.800 15.200 ;
        RECT 135.000 15.100 135.400 15.200 ;
        RECT 133.400 14.800 135.400 15.100 ;
        RECT 136.600 14.800 137.000 15.200 ;
        RECT 138.200 14.800 138.600 15.200 ;
        RECT 139.800 14.800 140.200 15.200 ;
        RECT 126.200 13.800 126.600 14.200 ;
        RECT 124.600 12.800 125.000 13.200 ;
        RECT 120.600 11.800 121.000 12.200 ;
        RECT 114.200 8.800 114.600 9.200 ;
        RECT 116.600 8.800 117.000 9.200 ;
        RECT 119.000 8.800 119.400 9.200 ;
        RECT 111.000 7.800 111.400 8.200 ;
        RECT 112.600 7.800 113.000 8.200 ;
        RECT 112.600 7.200 112.900 7.800 ;
        RECT 112.600 6.800 113.000 7.200 ;
        RECT 106.200 5.800 107.300 6.100 ;
        RECT 107.800 5.800 108.200 6.200 ;
        RECT 110.200 5.800 110.600 6.200 ;
        RECT 111.000 6.100 111.400 6.200 ;
        RECT 111.800 6.100 112.200 6.200 ;
        RECT 111.000 5.800 112.200 6.100 ;
        RECT 114.200 6.100 114.500 8.800 ;
        RECT 127.800 8.200 128.100 14.800 ;
        RECT 128.600 13.800 129.000 14.200 ;
        RECT 135.000 14.100 135.400 14.200 ;
        RECT 136.600 14.100 137.000 14.200 ;
        RECT 137.400 14.100 137.800 14.200 ;
        RECT 135.000 13.800 136.100 14.100 ;
        RECT 136.600 13.800 137.800 14.100 ;
        RECT 128.600 13.200 128.900 13.800 ;
        RECT 135.800 13.200 136.100 13.800 ;
        RECT 128.600 12.800 129.000 13.200 ;
        RECT 131.000 12.800 131.400 13.200 ;
        RECT 134.200 13.100 134.600 13.200 ;
        RECT 135.000 13.100 135.400 13.200 ;
        RECT 134.200 12.800 135.400 13.100 ;
        RECT 135.800 12.800 136.200 13.200 ;
        RECT 131.000 12.200 131.300 12.800 ;
        RECT 131.000 11.800 131.400 12.200 ;
        RECT 137.400 11.800 137.800 12.200 ;
        RECT 129.400 8.800 129.800 9.200 ;
        RECT 134.200 8.800 134.600 9.200 ;
        RECT 115.000 8.100 115.400 8.200 ;
        RECT 116.600 8.100 117.000 8.200 ;
        RECT 115.000 7.800 117.000 8.100 ;
        RECT 122.200 7.800 122.600 8.200 ;
        RECT 127.800 7.800 128.200 8.200 ;
        RECT 122.200 7.200 122.500 7.800 ;
        RECT 129.400 7.200 129.700 8.800 ;
        RECT 134.200 8.200 134.500 8.800 ;
        RECT 134.200 7.800 134.600 8.200 ;
        RECT 136.600 7.800 137.000 8.200 ;
        RECT 136.600 7.200 136.900 7.800 ;
        RECT 137.400 7.200 137.700 11.800 ;
        RECT 138.200 9.200 138.500 14.800 ;
        RECT 139.800 12.200 140.100 14.800 ;
        RECT 140.600 14.200 140.900 17.800 ;
        RECT 140.600 13.800 141.000 14.200 ;
        RECT 139.800 11.800 140.200 12.200 ;
        RECT 141.400 12.100 141.700 25.800 ;
        RECT 143.000 23.200 143.300 26.800 ;
        RECT 146.200 26.200 146.500 31.800 ;
        RECT 147.800 28.200 148.100 33.800 ;
        RECT 150.200 29.200 150.500 45.800 ;
        RECT 150.200 28.800 150.600 29.200 ;
        RECT 147.800 27.800 148.200 28.200 ;
        RECT 146.200 25.800 146.600 26.200 ;
        RECT 146.200 24.800 146.600 25.200 ;
        RECT 143.000 22.800 143.400 23.200 ;
        RECT 146.200 19.200 146.500 24.800 ;
        RECT 146.200 18.800 146.600 19.200 ;
        RECT 147.800 15.800 148.200 16.200 ;
        RECT 147.800 15.200 148.100 15.800 ;
        RECT 143.800 15.100 144.200 15.200 ;
        RECT 143.800 14.800 144.900 15.100 ;
        RECT 147.800 14.800 148.200 15.200 ;
        RECT 148.600 15.100 149.000 15.200 ;
        RECT 149.400 15.100 149.800 15.200 ;
        RECT 148.600 14.800 149.800 15.100 ;
        RECT 142.200 13.800 142.600 14.200 ;
        RECT 142.200 13.200 142.500 13.800 ;
        RECT 142.200 12.800 142.600 13.200 ;
        RECT 143.000 12.800 143.400 13.200 ;
        RECT 141.400 11.800 142.500 12.100 ;
        RECT 141.400 10.800 141.800 11.200 ;
        RECT 141.400 9.200 141.700 10.800 ;
        RECT 138.200 8.800 138.600 9.200 ;
        RECT 141.400 8.800 141.800 9.200 ;
        RECT 142.200 8.200 142.500 11.800 ;
        RECT 143.000 11.200 143.300 12.800 ;
        RECT 143.000 10.800 143.400 11.200 ;
        RECT 144.600 9.200 144.900 14.800 ;
        RECT 144.600 8.800 145.000 9.200 ;
        RECT 142.200 7.800 142.600 8.200 ;
        RECT 143.800 7.800 144.200 8.200 ;
        RECT 145.400 7.800 145.800 8.200 ;
        RECT 146.200 7.800 146.600 8.200 ;
        RECT 143.800 7.200 144.100 7.800 ;
        RECT 145.400 7.200 145.700 7.800 ;
        RECT 146.200 7.200 146.500 7.800 ;
        RECT 115.000 7.100 115.400 7.200 ;
        RECT 115.800 7.100 116.200 7.200 ;
        RECT 115.000 6.800 116.200 7.100 ;
        RECT 117.400 7.100 117.800 7.200 ;
        RECT 118.200 7.100 118.600 7.200 ;
        RECT 117.400 6.800 118.600 7.100 ;
        RECT 119.800 6.800 120.200 7.200 ;
        RECT 122.200 6.800 122.600 7.200 ;
        RECT 123.000 7.100 123.400 7.200 ;
        RECT 123.800 7.100 124.200 7.200 ;
        RECT 123.000 6.800 124.200 7.100 ;
        RECT 128.600 7.100 129.000 7.200 ;
        RECT 129.400 7.100 129.800 7.200 ;
        RECT 128.600 6.800 129.800 7.100 ;
        RECT 132.600 7.100 133.000 7.200 ;
        RECT 132.600 6.800 133.700 7.100 ;
        RECT 136.600 6.800 137.000 7.200 ;
        RECT 137.400 6.800 137.800 7.200 ;
        RECT 143.800 6.800 144.200 7.200 ;
        RECT 145.400 6.800 145.800 7.200 ;
        RECT 146.200 6.800 146.600 7.200 ;
        RECT 147.800 7.100 148.200 7.200 ;
        RECT 148.600 7.100 149.000 7.200 ;
        RECT 147.800 6.800 149.000 7.100 ;
        RECT 119.800 6.200 120.100 6.800 ;
        RECT 115.000 6.100 115.400 6.200 ;
        RECT 114.200 5.800 115.400 6.100 ;
        RECT 119.800 5.800 120.200 6.200 ;
        RECT 120.600 6.100 121.000 6.200 ;
        RECT 121.400 6.100 121.800 6.200 ;
        RECT 120.600 5.800 121.800 6.100 ;
        RECT 129.400 6.100 129.800 6.200 ;
        RECT 130.200 6.100 130.600 6.200 ;
        RECT 129.400 5.800 130.600 6.100 ;
        RECT 131.800 6.100 132.200 6.200 ;
        RECT 132.600 6.100 133.000 6.200 ;
        RECT 131.800 5.800 133.000 6.100 ;
        RECT 86.200 5.200 86.500 5.800 ;
        RECT 39.800 4.800 40.200 5.200 ;
        RECT 78.200 5.100 78.600 5.200 ;
        RECT 79.000 5.100 79.400 5.200 ;
        RECT 79.800 5.100 80.200 5.200 ;
        RECT 78.200 4.800 80.200 5.100 ;
        RECT 81.400 4.800 81.800 5.200 ;
        RECT 86.200 4.800 86.600 5.200 ;
        RECT 94.200 5.100 94.500 5.800 ;
        RECT 95.800 5.100 96.100 5.800 ;
        RECT 94.200 4.800 96.100 5.100 ;
        RECT 107.800 5.200 108.100 5.800 ;
        RECT 133.400 5.200 133.700 6.800 ;
        RECT 137.400 6.200 137.700 6.800 ;
        RECT 137.400 5.800 137.800 6.200 ;
        RECT 139.800 5.800 140.200 6.200 ;
        RECT 142.200 6.100 142.600 6.200 ;
        RECT 143.000 6.100 143.400 6.200 ;
        RECT 142.200 5.800 143.400 6.100 ;
        RECT 146.200 6.100 146.600 6.200 ;
        RECT 147.000 6.100 147.400 6.200 ;
        RECT 146.200 5.800 147.400 6.100 ;
        RECT 139.800 5.200 140.100 5.800 ;
        RECT 149.400 5.200 149.700 14.800 ;
        RECT 107.800 4.800 108.200 5.200 ;
        RECT 131.000 5.100 131.400 5.200 ;
        RECT 131.800 5.100 132.200 5.200 ;
        RECT 131.000 4.800 132.200 5.100 ;
        RECT 133.400 4.800 133.800 5.200 ;
        RECT 139.800 4.800 140.200 5.200 ;
        RECT 149.400 4.800 149.800 5.200 ;
      LAYER via2 ;
        RECT 20.600 126.800 21.000 127.200 ;
        RECT 11.800 125.800 12.200 126.200 ;
        RECT 20.600 125.800 21.000 126.200 ;
        RECT 13.400 124.800 13.800 125.200 ;
        RECT 12.600 123.800 13.000 124.200 ;
        RECT 19.000 121.800 19.400 122.200 ;
        RECT 23.000 123.800 23.400 124.200 ;
        RECT 2.200 116.800 2.600 117.200 ;
        RECT 12.600 115.800 13.000 116.200 ;
        RECT 4.600 114.800 5.000 115.200 ;
        RECT 3.800 105.800 4.200 106.200 ;
        RECT 1.400 104.800 1.800 105.200 ;
        RECT 7.800 98.800 8.200 99.200 ;
        RECT 14.200 106.800 14.600 107.200 ;
        RECT 16.600 106.800 17.000 107.200 ;
        RECT 2.200 96.800 2.600 97.200 ;
        RECT 9.400 95.800 9.800 96.200 ;
        RECT 25.400 123.800 25.800 124.200 ;
        RECT 31.000 125.800 31.400 126.200 ;
        RECT 35.800 125.800 36.200 126.200 ;
        RECT 63.800 126.800 64.200 127.200 ;
        RECT 67.000 126.800 67.400 127.200 ;
        RECT 40.600 108.800 41.000 109.200 ;
        RECT 31.800 103.800 32.200 104.200 ;
        RECT 43.000 104.800 43.400 105.200 ;
        RECT 58.200 113.800 58.600 114.200 ;
        RECT 60.600 113.800 61.000 114.200 ;
        RECT 64.600 113.800 65.000 114.200 ;
        RECT 47.800 103.800 48.200 104.200 ;
        RECT 58.200 105.800 58.600 106.200 ;
        RECT 51.800 98.800 52.200 99.200 ;
        RECT 7.000 86.800 7.400 87.200 ;
        RECT 10.200 75.800 10.600 76.200 ;
        RECT 39.800 96.800 40.200 97.200 ;
        RECT 12.600 86.800 13.000 87.200 ;
        RECT 25.400 86.800 25.800 87.200 ;
        RECT 19.000 83.800 19.400 84.200 ;
        RECT 39.000 94.800 39.400 95.200 ;
        RECT 42.200 93.800 42.600 94.200 ;
        RECT 33.400 91.800 33.800 92.200 ;
        RECT 37.400 88.800 37.800 89.200 ;
        RECT 34.200 86.800 34.600 87.200 ;
        RECT 17.400 75.800 17.800 76.200 ;
        RECT 25.400 75.800 25.800 76.200 ;
        RECT 20.600 74.800 21.000 75.200 ;
        RECT 8.600 66.800 9.000 67.200 ;
        RECT 4.600 56.800 5.000 57.200 ;
        RECT 3.800 54.800 4.200 55.200 ;
        RECT 24.600 67.800 25.000 68.200 ;
        RECT 38.200 86.800 38.600 87.200 ;
        RECT 39.800 86.800 40.200 87.200 ;
        RECT 48.600 86.800 49.000 87.200 ;
        RECT 53.400 86.800 53.800 87.200 ;
        RECT 31.800 84.800 32.200 85.200 ;
        RECT 43.800 84.800 44.200 85.200 ;
        RECT 35.800 83.800 36.200 84.200 ;
        RECT 39.000 73.800 39.400 74.200 ;
        RECT 62.200 94.800 62.600 95.200 ;
        RECT 59.000 87.800 59.400 88.200 ;
        RECT 69.400 106.800 69.800 107.200 ;
        RECT 99.800 121.800 100.200 122.200 ;
        RECT 121.400 127.800 121.800 128.200 ;
        RECT 107.000 118.800 107.400 119.200 ;
        RECT 112.600 115.800 113.000 116.200 ;
        RECT 121.400 115.800 121.800 116.200 ;
        RECT 119.800 113.800 120.200 114.200 ;
        RECT 73.400 107.800 73.800 108.200 ;
        RECT 91.000 107.800 91.400 108.200 ;
        RECT 73.400 106.800 73.800 107.200 ;
        RECT 67.000 104.800 67.400 105.200 ;
        RECT 72.600 104.800 73.000 105.200 ;
        RECT 71.000 96.800 71.400 97.200 ;
        RECT 91.800 105.800 92.200 106.200 ;
        RECT 85.400 103.800 85.800 104.200 ;
        RECT 86.200 98.800 86.600 99.200 ;
        RECT 39.800 70.800 40.200 71.200 ;
        RECT 19.800 65.800 20.200 66.200 ;
        RECT 39.800 64.800 40.200 65.200 ;
        RECT 6.200 44.800 6.600 45.200 ;
        RECT 3.000 34.800 3.400 35.200 ;
        RECT 4.600 34.800 5.000 35.200 ;
        RECT 8.600 34.800 9.000 35.200 ;
        RECT 3.800 33.800 4.200 34.200 ;
        RECT 26.200 62.800 26.600 63.200 ;
        RECT 23.000 56.800 23.400 57.200 ;
        RECT 15.000 53.800 15.400 54.200 ;
        RECT 36.600 56.800 37.000 57.200 ;
        RECT 17.400 45.800 17.800 46.200 ;
        RECT 28.600 52.800 29.000 53.200 ;
        RECT 35.800 54.800 36.200 55.200 ;
        RECT 43.800 47.800 44.200 48.200 ;
        RECT 31.000 46.800 31.400 47.200 ;
        RECT 30.200 45.800 30.600 46.200 ;
        RECT 17.400 32.800 17.800 33.200 ;
        RECT 21.400 34.800 21.800 35.200 ;
        RECT 25.400 35.800 25.800 36.200 ;
        RECT 43.800 46.800 44.200 47.200 ;
        RECT 79.000 96.800 79.400 97.200 ;
        RECT 75.800 94.800 76.200 95.200 ;
        RECT 80.600 94.800 81.000 95.200 ;
        RECT 72.600 92.800 73.000 93.200 ;
        RECT 78.200 93.800 78.600 94.200 ;
        RECT 68.600 76.800 69.000 77.200 ;
        RECT 121.400 107.800 121.800 108.200 ;
        RECT 119.800 101.800 120.200 102.200 ;
        RECT 92.600 93.800 93.000 94.200 ;
        RECT 74.200 88.800 74.600 89.200 ;
        RECT 93.400 88.800 93.800 89.200 ;
        RECT 64.600 67.800 65.000 68.200 ;
        RECT 70.200 67.800 70.600 68.200 ;
        RECT 63.800 65.800 64.200 66.200 ;
        RECT 58.200 58.800 58.600 59.200 ;
        RECT 60.600 54.800 61.000 55.200 ;
        RECT 58.200 46.800 58.600 47.200 ;
        RECT 61.400 46.800 61.800 47.200 ;
        RECT 46.200 45.800 46.600 46.200 ;
        RECT 32.600 32.800 33.000 33.200 ;
        RECT 30.200 26.800 30.600 27.200 ;
        RECT 19.800 23.800 20.200 24.200 ;
        RECT 6.200 14.800 6.600 15.200 ;
        RECT 14.200 15.800 14.600 16.200 ;
        RECT 13.400 14.800 13.800 15.200 ;
        RECT 15.800 5.800 16.200 6.200 ;
        RECT 37.400 21.800 37.800 22.200 ;
        RECT 29.400 14.800 29.800 15.200 ;
        RECT 36.600 16.800 37.000 17.200 ;
        RECT 30.200 13.800 30.600 14.200 ;
        RECT 106.200 86.800 106.600 87.200 ;
        RECT 119.800 93.800 120.200 94.200 ;
        RECT 123.800 106.800 124.200 107.200 ;
        RECT 139.800 113.800 140.200 114.200 ;
        RECT 141.400 112.800 141.800 113.200 ;
        RECT 142.200 105.800 142.600 106.200 ;
        RECT 122.200 92.800 122.600 93.200 ;
        RECT 118.200 87.800 118.600 88.200 ;
        RECT 117.400 85.800 117.800 86.200 ;
        RECT 81.400 55.800 81.800 56.200 ;
        RECT 76.600 51.800 77.000 52.200 ;
        RECT 93.400 61.800 93.800 62.200 ;
        RECT 81.400 46.800 81.800 47.200 ;
        RECT 71.000 34.800 71.400 35.200 ;
        RECT 97.400 54.800 97.800 55.200 ;
        RECT 91.800 45.800 92.200 46.200 ;
        RECT 111.800 72.800 112.200 73.200 ;
        RECT 115.000 69.800 115.400 70.200 ;
        RECT 115.800 67.800 116.200 68.200 ;
        RECT 147.000 94.800 147.400 95.200 ;
        RECT 130.200 73.800 130.600 74.200 ;
        RECT 123.000 67.800 123.400 68.200 ;
        RECT 127.800 65.800 128.200 66.200 ;
        RECT 124.600 64.800 125.000 65.200 ;
        RECT 119.000 55.800 119.400 56.200 ;
        RECT 137.400 53.800 137.800 54.200 ;
        RECT 94.200 44.800 94.600 45.200 ;
        RECT 55.800 24.800 56.200 25.200 ;
        RECT 38.200 13.800 38.600 14.200 ;
        RECT 46.200 13.800 46.600 14.200 ;
        RECT 26.200 4.800 26.600 5.200 ;
        RECT 45.400 6.800 45.800 7.200 ;
        RECT 31.000 4.800 31.400 5.200 ;
        RECT 67.000 25.800 67.400 26.200 ;
        RECT 84.600 32.800 85.000 33.200 ;
        RECT 107.800 35.800 108.200 36.200 ;
        RECT 121.400 46.800 121.800 47.200 ;
        RECT 122.200 45.800 122.600 46.200 ;
        RECT 145.400 54.800 145.800 55.200 ;
        RECT 147.000 54.800 147.400 55.200 ;
        RECT 143.000 53.800 143.400 54.200 ;
        RECT 135.000 46.800 135.400 47.200 ;
        RECT 119.800 34.800 120.200 35.200 ;
        RECT 115.800 27.800 116.200 28.200 ;
        RECT 98.200 26.800 98.600 27.200 ;
        RECT 100.600 26.800 101.000 27.200 ;
        RECT 75.000 16.800 75.400 17.200 ;
        RECT 69.400 11.800 69.800 12.200 ;
        RECT 77.400 15.800 77.800 16.200 ;
        RECT 70.200 7.800 70.600 8.200 ;
        RECT 54.200 6.800 54.600 7.200 ;
        RECT 79.800 6.800 80.200 7.200 ;
        RECT 37.400 5.800 37.800 6.200 ;
        RECT 48.600 5.800 49.000 6.200 ;
        RECT 71.000 5.800 71.400 6.200 ;
        RECT 74.200 5.800 74.600 6.200 ;
        RECT 96.600 8.800 97.000 9.200 ;
        RECT 103.000 26.600 103.400 27.000 ;
        RECT 119.000 26.800 119.400 27.200 ;
        RECT 138.200 35.800 138.600 36.200 ;
        RECT 133.400 32.800 133.800 33.200 ;
        RECT 124.600 25.800 125.000 26.200 ;
        RECT 106.200 16.800 106.600 17.200 ;
        RECT 107.000 15.800 107.400 16.200 ;
        RECT 110.200 13.800 110.600 14.200 ;
        RECT 102.200 5.800 102.600 6.200 ;
        RECT 103.800 5.800 104.200 6.200 ;
        RECT 119.800 24.800 120.200 25.200 ;
        RECT 128.600 16.800 129.000 17.200 ;
        RECT 140.600 33.800 141.000 34.200 ;
        RECT 150.200 50.800 150.600 51.200 ;
        RECT 142.200 26.800 142.600 27.200 ;
        RECT 139.000 15.800 139.400 16.200 ;
        RECT 149.400 14.800 149.800 15.200 ;
        RECT 118.200 6.800 118.600 7.200 ;
        RECT 123.800 6.800 124.200 7.200 ;
        RECT 148.600 6.800 149.000 7.200 ;
        RECT 79.000 4.800 79.400 5.200 ;
      LAYER metal3 ;
        RECT 10.200 129.100 10.600 129.200 ;
        RECT 46.200 129.100 46.600 129.200 ;
        RECT 10.200 128.800 46.600 129.100 ;
        RECT 7.000 127.800 7.400 128.200 ;
        RECT 13.400 128.100 13.800 128.200 ;
        RECT 23.800 128.100 24.200 128.200 ;
        RECT 27.000 128.100 27.400 128.200 ;
        RECT 13.400 127.800 20.100 128.100 ;
        RECT 23.800 127.800 27.400 128.100 ;
        RECT 27.800 127.800 28.200 128.200 ;
        RECT 39.800 128.100 40.200 128.200 ;
        RECT 40.600 128.100 41.000 128.200 ;
        RECT 39.800 127.800 41.000 128.100 ;
        RECT 41.400 128.100 41.800 128.200 ;
        RECT 56.600 128.100 57.000 128.200 ;
        RECT 41.400 127.800 57.000 128.100 ;
        RECT 62.200 128.100 62.600 128.200 ;
        RECT 65.400 128.100 65.800 128.200 ;
        RECT 62.200 127.800 65.800 128.100 ;
        RECT 121.400 128.100 121.800 128.200 ;
        RECT 137.400 128.100 137.800 128.200 ;
        RECT 121.400 127.800 137.800 128.100 ;
        RECT 0.600 126.800 1.000 127.200 ;
        RECT 1.400 127.100 1.800 127.200 ;
        RECT 3.800 127.100 4.200 127.200 ;
        RECT 1.400 126.800 4.200 127.100 ;
        RECT 7.000 127.100 7.300 127.800 ;
        RECT 14.200 127.100 14.600 127.200 ;
        RECT 7.000 126.800 14.600 127.100 ;
        RECT 15.000 127.100 15.400 127.200 ;
        RECT 18.200 127.100 18.600 127.200 ;
        RECT 15.000 126.800 18.600 127.100 ;
        RECT 19.800 127.100 20.100 127.800 ;
        RECT 20.600 127.100 21.000 127.200 ;
        RECT 27.800 127.100 28.100 127.800 ;
        RECT 19.800 126.800 28.100 127.100 ;
        RECT 31.800 127.100 32.200 127.200 ;
        RECT 41.400 127.100 41.800 127.200 ;
        RECT 31.800 126.800 41.800 127.100 ;
        RECT 45.400 127.100 45.800 127.200 ;
        RECT 51.000 127.100 51.400 127.200 ;
        RECT 45.400 126.800 51.400 127.100 ;
        RECT 59.800 127.100 60.200 127.200 ;
        RECT 63.800 127.100 64.200 127.200 ;
        RECT 59.800 126.800 64.200 127.100 ;
        RECT 64.600 127.100 65.000 127.200 ;
        RECT 65.400 127.100 65.800 127.200 ;
        RECT 64.600 126.800 65.800 127.100 ;
        RECT 67.000 127.100 67.400 127.200 ;
        RECT 68.600 127.100 69.000 127.200 ;
        RECT 67.000 126.800 69.000 127.100 ;
        RECT 73.400 127.100 73.800 127.200 ;
        RECT 74.200 127.100 74.600 127.200 ;
        RECT 73.400 126.800 74.600 127.100 ;
        RECT 77.400 127.100 77.800 127.200 ;
        RECT 84.600 127.100 85.000 127.200 ;
        RECT 77.400 126.800 85.000 127.100 ;
        RECT 89.400 126.800 89.800 127.200 ;
        RECT 0.600 126.100 0.900 126.800 ;
        RECT 89.400 126.200 89.700 126.800 ;
        RECT 9.400 126.100 9.800 126.200 ;
        RECT 11.800 126.100 12.200 126.200 ;
        RECT 0.600 125.800 12.200 126.100 ;
        RECT 15.800 126.100 16.200 126.200 ;
        RECT 20.600 126.100 21.000 126.200 ;
        RECT 31.000 126.100 31.400 126.200 ;
        RECT 35.800 126.100 36.200 126.200 ;
        RECT 39.800 126.100 40.200 126.200 ;
        RECT 42.200 126.100 42.600 126.200 ;
        RECT 15.800 125.800 30.500 126.100 ;
        RECT 31.000 125.800 42.600 126.100 ;
        RECT 45.400 126.100 45.800 126.200 ;
        RECT 50.200 126.100 50.600 126.200 ;
        RECT 45.400 125.800 50.600 126.100 ;
        RECT 61.400 126.100 61.800 126.200 ;
        RECT 65.400 126.100 65.800 126.200 ;
        RECT 71.800 126.100 72.200 126.200 ;
        RECT 75.800 126.100 76.200 126.200 ;
        RECT 80.600 126.100 81.000 126.200 ;
        RECT 61.400 125.800 81.000 126.100 ;
        RECT 89.400 125.800 89.800 126.200 ;
        RECT 95.000 126.100 95.400 126.200 ;
        RECT 103.000 126.100 103.400 126.200 ;
        RECT 122.200 126.100 122.600 126.200 ;
        RECT 95.000 125.800 122.600 126.100 ;
        RECT 8.600 125.100 9.000 125.200 ;
        RECT 9.400 125.100 9.800 125.200 ;
        RECT 13.400 125.100 13.800 125.200 ;
        RECT 17.400 125.100 17.800 125.200 ;
        RECT 8.600 124.800 9.800 125.100 ;
        RECT 12.600 124.800 17.800 125.100 ;
        RECT 23.800 125.100 24.200 125.200 ;
        RECT 26.200 125.100 26.600 125.200 ;
        RECT 23.800 124.800 26.600 125.100 ;
        RECT 30.200 125.100 30.500 125.800 ;
        RECT 38.200 125.100 38.600 125.200 ;
        RECT 55.000 125.100 55.400 125.200 ;
        RECT 30.200 124.800 55.400 125.100 ;
        RECT 55.800 125.100 56.200 125.200 ;
        RECT 73.400 125.100 73.800 125.200 ;
        RECT 81.400 125.100 81.800 125.200 ;
        RECT 87.000 125.100 87.400 125.200 ;
        RECT 55.800 124.800 87.400 125.100 ;
        RECT 103.000 125.100 103.400 125.200 ;
        RECT 143.800 125.100 144.200 125.200 ;
        RECT 103.000 124.800 144.200 125.100 ;
        RECT 147.800 124.800 148.200 125.200 ;
        RECT 147.800 124.200 148.100 124.800 ;
        RECT 2.200 124.100 2.600 124.200 ;
        RECT 3.800 124.100 4.200 124.200 ;
        RECT 9.400 124.100 9.800 124.200 ;
        RECT 2.200 123.800 9.800 124.100 ;
        RECT 12.600 124.100 13.000 124.200 ;
        RECT 23.000 124.100 23.400 124.200 ;
        RECT 12.600 123.800 23.400 124.100 ;
        RECT 25.400 124.100 25.800 124.200 ;
        RECT 36.600 124.100 37.000 124.200 ;
        RECT 25.400 123.800 37.000 124.100 ;
        RECT 38.200 124.100 38.600 124.200 ;
        RECT 40.600 124.100 41.000 124.200 ;
        RECT 38.200 123.800 41.000 124.100 ;
        RECT 41.400 124.100 41.800 124.200 ;
        RECT 42.200 124.100 42.600 124.200 ;
        RECT 41.400 123.800 42.600 124.100 ;
        RECT 47.800 124.100 48.200 124.200 ;
        RECT 51.000 124.100 51.400 124.200 ;
        RECT 72.600 124.100 73.000 124.200 ;
        RECT 47.800 123.800 73.000 124.100 ;
        RECT 147.800 123.800 148.200 124.200 ;
        RECT 70.200 123.200 70.500 123.800 ;
        RECT 17.400 123.100 17.800 123.200 ;
        RECT 27.000 123.100 27.400 123.200 ;
        RECT 17.400 122.800 27.400 123.100 ;
        RECT 29.400 123.100 29.800 123.200 ;
        RECT 35.800 123.100 36.200 123.200 ;
        RECT 44.600 123.100 45.000 123.200 ;
        RECT 59.800 123.100 60.200 123.200 ;
        RECT 29.400 122.800 60.200 123.100 ;
        RECT 70.200 122.800 70.600 123.200 ;
        RECT 19.000 122.100 19.400 122.200 ;
        RECT 32.600 122.100 33.000 122.200 ;
        RECT 19.000 121.800 33.000 122.100 ;
        RECT 99.800 122.100 100.200 122.200 ;
        RECT 141.400 122.100 141.800 122.200 ;
        RECT 99.800 121.800 141.800 122.100 ;
        RECT 3.000 121.100 3.400 121.200 ;
        RECT 6.200 121.100 6.600 121.200 ;
        RECT 38.200 121.100 38.600 121.200 ;
        RECT 3.000 120.800 38.600 121.100 ;
        RECT 55.000 121.100 55.400 121.200 ;
        RECT 112.600 121.100 113.000 121.200 ;
        RECT 55.000 120.800 113.000 121.100 ;
        RECT 113.400 121.100 113.800 121.200 ;
        RECT 118.200 121.100 118.600 121.200 ;
        RECT 140.600 121.100 141.000 121.200 ;
        RECT 113.400 120.800 141.000 121.100 ;
        RECT 55.000 120.100 55.400 120.200 ;
        RECT 59.800 120.100 60.200 120.200 ;
        RECT 55.000 119.800 60.200 120.100 ;
        RECT 64.600 120.100 65.000 120.200 ;
        RECT 79.000 120.100 79.400 120.200 ;
        RECT 64.600 119.800 79.400 120.100 ;
        RECT 116.600 120.100 117.000 120.200 ;
        RECT 127.800 120.100 128.200 120.200 ;
        RECT 116.600 119.800 128.200 120.100 ;
        RECT 19.800 119.100 20.200 119.200 ;
        RECT 55.800 119.100 56.200 119.200 ;
        RECT 67.800 119.100 68.200 119.200 ;
        RECT 19.800 118.800 56.200 119.100 ;
        RECT 59.000 118.800 68.200 119.100 ;
        RECT 74.200 119.100 74.600 119.200 ;
        RECT 105.400 119.100 105.800 119.200 ;
        RECT 74.200 118.800 105.800 119.100 ;
        RECT 107.000 119.100 107.400 119.200 ;
        RECT 108.600 119.100 109.000 119.200 ;
        RECT 107.000 118.800 109.000 119.100 ;
        RECT 59.000 118.200 59.300 118.800 ;
        RECT 7.000 118.100 7.400 118.200 ;
        RECT 23.800 118.100 24.200 118.200 ;
        RECT 7.000 117.800 24.200 118.100 ;
        RECT 27.000 117.800 27.400 118.200 ;
        RECT 34.200 118.100 34.600 118.200 ;
        RECT 39.000 118.100 39.400 118.200 ;
        RECT 42.200 118.100 42.600 118.200 ;
        RECT 59.000 118.100 59.400 118.200 ;
        RECT 34.200 117.800 59.400 118.100 ;
        RECT 71.800 117.800 72.200 118.200 ;
        RECT 81.400 118.100 81.800 118.200 ;
        RECT 120.600 118.100 121.000 118.200 ;
        RECT 81.400 117.800 121.000 118.100 ;
        RECT 2.200 117.100 2.600 117.200 ;
        RECT 3.800 117.100 4.200 117.200 ;
        RECT 4.600 117.100 5.000 117.200 ;
        RECT 2.200 116.800 5.000 117.100 ;
        RECT 11.800 117.100 12.200 117.200 ;
        RECT 15.000 117.100 15.400 117.200 ;
        RECT 11.800 116.800 15.400 117.100 ;
        RECT 16.600 117.100 17.000 117.200 ;
        RECT 27.000 117.100 27.300 117.800 ;
        RECT 36.600 117.100 37.000 117.200 ;
        RECT 43.000 117.100 43.400 117.200 ;
        RECT 16.600 116.800 25.700 117.100 ;
        RECT 27.000 116.800 43.400 117.100 ;
        RECT 71.800 117.100 72.100 117.800 ;
        RECT 74.200 117.100 74.600 117.200 ;
        RECT 71.800 116.800 74.600 117.100 ;
        RECT 101.400 117.100 101.800 117.200 ;
        RECT 109.400 117.100 109.800 117.200 ;
        RECT 101.400 116.800 109.800 117.100 ;
        RECT 25.400 116.200 25.700 116.800 ;
        RECT 6.200 116.100 6.600 116.200 ;
        RECT 11.000 116.100 11.400 116.200 ;
        RECT 6.200 115.800 11.400 116.100 ;
        RECT 12.600 116.100 13.000 116.200 ;
        RECT 14.200 116.100 14.600 116.200 ;
        RECT 12.600 115.800 14.600 116.100 ;
        RECT 20.600 116.100 21.000 116.200 ;
        RECT 22.200 116.100 22.600 116.200 ;
        RECT 20.600 115.800 22.600 116.100 ;
        RECT 25.400 115.800 25.800 116.200 ;
        RECT 30.200 116.100 30.600 116.200 ;
        RECT 33.400 116.100 33.800 116.200 ;
        RECT 30.200 115.800 33.800 116.100 ;
        RECT 63.000 116.100 63.400 116.200 ;
        RECT 67.000 116.100 67.400 116.200 ;
        RECT 63.000 115.800 67.400 116.100 ;
        RECT 108.600 116.100 109.000 116.200 ;
        RECT 111.000 116.100 111.400 116.200 ;
        RECT 108.600 115.800 111.400 116.100 ;
        RECT 112.600 116.100 113.000 116.200 ;
        RECT 114.200 116.100 114.600 116.200 ;
        RECT 119.800 116.100 120.200 116.200 ;
        RECT 112.600 115.800 120.200 116.100 ;
        RECT 121.400 116.100 121.800 116.200 ;
        RECT 128.600 116.100 129.000 116.200 ;
        RECT 121.400 115.800 129.000 116.100 ;
        RECT 2.200 114.800 2.600 115.200 ;
        RECT 4.600 115.100 5.000 115.200 ;
        RECT 7.000 115.100 7.400 115.200 ;
        RECT 15.000 115.100 15.400 115.200 ;
        RECT 23.800 115.100 24.200 115.200 ;
        RECT 4.600 114.800 24.200 115.100 ;
        RECT 33.400 115.100 33.800 115.200 ;
        RECT 35.800 115.100 36.200 115.200 ;
        RECT 42.200 115.100 42.600 115.200 ;
        RECT 33.400 114.800 42.600 115.100 ;
        RECT 61.400 115.100 61.800 115.200 ;
        RECT 66.200 115.100 66.600 115.200 ;
        RECT 61.400 114.800 66.600 115.100 ;
        RECT 67.000 115.100 67.400 115.200 ;
        RECT 67.800 115.100 68.200 115.200 ;
        RECT 67.000 114.800 68.200 115.100 ;
        RECT 70.200 115.100 70.600 115.200 ;
        RECT 75.000 115.100 75.400 115.200 ;
        RECT 77.400 115.100 77.800 115.200 ;
        RECT 70.200 114.800 77.800 115.100 ;
        RECT 104.600 115.100 105.000 115.200 ;
        RECT 109.400 115.100 109.800 115.200 ;
        RECT 104.600 114.800 109.800 115.100 ;
        RECT 112.600 115.100 113.000 115.200 ;
        RECT 116.600 115.100 117.000 115.200 ;
        RECT 112.600 114.800 117.000 115.100 ;
        RECT 117.400 115.100 117.800 115.200 ;
        RECT 119.800 115.100 120.200 115.200 ;
        RECT 117.400 114.800 120.200 115.100 ;
        RECT 120.600 114.800 121.000 115.200 ;
        RECT 2.200 114.200 2.500 114.800 ;
        RECT 120.600 114.200 120.900 114.800 ;
        RECT 2.200 113.800 2.600 114.200 ;
        RECT 3.000 114.100 3.400 114.200 ;
        RECT 16.600 114.100 17.000 114.200 ;
        RECT 28.600 114.100 29.000 114.200 ;
        RECT 3.000 113.800 17.000 114.100 ;
        RECT 21.400 113.800 29.000 114.100 ;
        RECT 31.800 114.100 32.200 114.200 ;
        RECT 40.600 114.100 41.000 114.200 ;
        RECT 31.800 113.800 41.000 114.100 ;
        RECT 58.200 114.100 58.600 114.200 ;
        RECT 60.600 114.100 61.000 114.200 ;
        RECT 58.200 113.800 61.000 114.100 ;
        RECT 63.000 113.800 63.400 114.200 ;
        RECT 64.600 114.100 65.000 114.200 ;
        RECT 67.800 114.100 68.200 114.200 ;
        RECT 73.400 114.100 73.800 114.200 ;
        RECT 64.600 113.800 73.800 114.100 ;
        RECT 104.600 114.100 105.000 114.200 ;
        RECT 107.000 114.100 107.400 114.200 ;
        RECT 114.200 114.100 114.600 114.200 ;
        RECT 119.800 114.100 120.200 114.200 ;
        RECT 104.600 113.800 120.200 114.100 ;
        RECT 120.600 113.800 121.000 114.200 ;
        RECT 139.800 114.100 140.200 114.200 ;
        RECT 140.600 114.100 141.000 114.200 ;
        RECT 139.800 113.800 141.000 114.100 ;
        RECT 21.400 113.200 21.700 113.800 ;
        RECT 2.200 113.100 2.600 113.200 ;
        RECT 5.400 113.100 5.800 113.200 ;
        RECT 2.200 112.800 5.800 113.100 ;
        RECT 11.000 113.100 11.400 113.200 ;
        RECT 17.400 113.100 17.800 113.200 ;
        RECT 11.000 112.800 17.800 113.100 ;
        RECT 21.400 112.800 21.800 113.200 ;
        RECT 23.800 113.100 24.200 113.200 ;
        RECT 29.400 113.100 29.800 113.200 ;
        RECT 34.200 113.100 34.600 113.200 ;
        RECT 23.800 112.800 34.600 113.100 ;
        RECT 36.600 113.100 37.000 113.200 ;
        RECT 39.800 113.100 40.200 113.200 ;
        RECT 36.600 112.800 40.200 113.100 ;
        RECT 54.200 113.100 54.600 113.200 ;
        RECT 55.800 113.100 56.200 113.200 ;
        RECT 54.200 112.800 56.200 113.100 ;
        RECT 63.000 113.100 63.300 113.800 ;
        RECT 63.800 113.100 64.200 113.200 ;
        RECT 63.000 112.800 64.200 113.100 ;
        RECT 66.200 113.100 66.600 113.200 ;
        RECT 69.400 113.100 69.800 113.200 ;
        RECT 83.800 113.100 84.200 113.200 ;
        RECT 66.200 112.800 84.200 113.100 ;
        RECT 98.200 113.100 98.600 113.200 ;
        RECT 102.200 113.100 102.600 113.200 ;
        RECT 98.200 112.800 102.600 113.100 ;
        RECT 118.200 113.100 118.600 113.200 ;
        RECT 139.800 113.100 140.200 113.200 ;
        RECT 118.200 112.800 140.200 113.100 ;
        RECT 141.400 113.100 141.800 113.200 ;
        RECT 143.800 113.100 144.200 113.200 ;
        RECT 141.400 112.800 144.200 113.100 ;
        RECT 19.000 112.100 19.400 112.200 ;
        RECT 30.200 112.100 30.600 112.200 ;
        RECT 19.000 111.800 30.600 112.100 ;
        RECT 34.200 112.100 34.600 112.200 ;
        RECT 43.000 112.100 43.400 112.200 ;
        RECT 34.200 111.800 43.400 112.100 ;
        RECT 45.400 112.100 45.800 112.200 ;
        RECT 55.800 112.100 56.200 112.200 ;
        RECT 45.400 111.800 56.200 112.100 ;
        RECT 59.800 112.100 60.200 112.200 ;
        RECT 71.000 112.100 71.400 112.200 ;
        RECT 80.600 112.100 81.000 112.200 ;
        RECT 59.800 111.800 81.000 112.100 ;
        RECT 95.800 112.100 96.200 112.200 ;
        RECT 99.800 112.100 100.200 112.200 ;
        RECT 95.800 111.800 100.200 112.100 ;
        RECT 20.600 111.100 21.000 111.200 ;
        RECT 27.000 111.100 27.400 111.200 ;
        RECT 20.600 110.800 27.400 111.100 ;
        RECT 31.800 111.100 32.200 111.200 ;
        RECT 35.000 111.100 35.400 111.200 ;
        RECT 56.600 111.100 57.000 111.200 ;
        RECT 31.800 110.800 57.000 111.100 ;
        RECT 81.400 111.100 81.800 111.200 ;
        RECT 87.000 111.100 87.400 111.200 ;
        RECT 81.400 110.800 87.400 111.100 ;
        RECT 89.400 111.100 89.800 111.200 ;
        RECT 92.600 111.100 93.000 111.200 ;
        RECT 89.400 110.800 93.000 111.100 ;
        RECT 147.000 110.800 147.400 111.200 ;
        RECT 23.000 110.100 23.400 110.200 ;
        RECT 31.800 110.100 32.100 110.800 ;
        RECT 147.000 110.200 147.300 110.800 ;
        RECT 23.000 109.800 32.100 110.100 ;
        RECT 32.600 110.100 33.000 110.200 ;
        RECT 91.800 110.100 92.200 110.200 ;
        RECT 32.600 109.800 92.200 110.100 ;
        RECT 111.000 110.100 111.400 110.200 ;
        RECT 145.400 110.100 145.800 110.200 ;
        RECT 111.000 109.800 145.800 110.100 ;
        RECT 147.000 109.800 147.400 110.200 ;
        RECT 8.600 109.100 9.000 109.200 ;
        RECT 11.000 109.100 11.400 109.200 ;
        RECT 25.400 109.100 25.800 109.200 ;
        RECT 40.600 109.100 41.000 109.200 ;
        RECT 8.600 108.800 16.900 109.100 ;
        RECT 25.400 108.800 41.000 109.100 ;
        RECT 51.800 109.100 52.200 109.200 ;
        RECT 60.600 109.100 61.000 109.200 ;
        RECT 51.800 108.800 61.000 109.100 ;
        RECT 62.200 109.100 62.600 109.200 ;
        RECT 76.600 109.100 77.000 109.200 ;
        RECT 86.200 109.100 86.600 109.200 ;
        RECT 62.200 108.800 66.500 109.100 ;
        RECT 76.600 108.800 100.100 109.100 ;
        RECT 16.600 108.200 16.900 108.800 ;
        RECT 66.200 108.200 66.500 108.800 ;
        RECT 99.800 108.200 100.100 108.800 ;
        RECT 5.400 108.100 5.800 108.200 ;
        RECT 12.600 108.100 13.000 108.200 ;
        RECT 5.400 107.800 13.000 108.100 ;
        RECT 16.600 107.800 17.000 108.200 ;
        RECT 19.800 108.100 20.200 108.200 ;
        RECT 25.400 108.100 25.800 108.200 ;
        RECT 19.800 107.800 25.800 108.100 ;
        RECT 28.600 108.100 29.000 108.200 ;
        RECT 35.000 108.100 35.400 108.200 ;
        RECT 28.600 107.800 35.400 108.100 ;
        RECT 51.000 108.100 51.400 108.200 ;
        RECT 55.000 108.100 55.400 108.200 ;
        RECT 64.600 108.100 65.000 108.200 ;
        RECT 51.000 107.800 65.000 108.100 ;
        RECT 66.200 107.800 66.600 108.200 ;
        RECT 71.000 108.100 71.400 108.200 ;
        RECT 73.400 108.100 73.800 108.200 ;
        RECT 91.000 108.100 91.400 108.200 ;
        RECT 96.600 108.100 97.000 108.200 ;
        RECT 71.000 107.800 78.500 108.100 ;
        RECT 91.000 107.800 97.000 108.100 ;
        RECT 99.800 107.800 100.200 108.200 ;
        RECT 121.400 108.100 121.800 108.200 ;
        RECT 130.200 108.100 130.600 108.200 ;
        RECT 121.400 107.800 130.600 108.100 ;
        RECT 78.200 107.200 78.500 107.800 ;
        RECT 3.800 107.100 4.200 107.200 ;
        RECT 8.600 107.100 9.000 107.200 ;
        RECT 14.200 107.100 14.600 107.200 ;
        RECT 15.800 107.100 16.200 107.200 ;
        RECT 16.600 107.100 17.000 107.200 ;
        RECT 3.800 106.800 17.000 107.100 ;
        RECT 24.600 107.100 25.000 107.200 ;
        RECT 32.600 107.100 33.000 107.200 ;
        RECT 24.600 106.800 33.000 107.100 ;
        RECT 34.200 107.100 34.600 107.200 ;
        RECT 39.000 107.100 39.400 107.200 ;
        RECT 43.800 107.100 44.200 107.200 ;
        RECT 46.200 107.100 46.600 107.200 ;
        RECT 34.200 106.800 46.600 107.100 ;
        RECT 47.000 107.100 47.400 107.200 ;
        RECT 51.000 107.100 51.400 107.200 ;
        RECT 47.000 106.800 51.400 107.100 ;
        RECT 55.800 107.100 56.200 107.200 ;
        RECT 58.200 107.100 58.600 107.200 ;
        RECT 55.800 106.800 58.600 107.100 ;
        RECT 67.800 106.800 68.200 107.200 ;
        RECT 69.400 107.100 69.800 107.200 ;
        RECT 71.800 107.100 72.200 107.200 ;
        RECT 73.400 107.100 73.800 107.200 ;
        RECT 69.400 106.800 73.800 107.100 ;
        RECT 78.200 106.800 78.600 107.200 ;
        RECT 87.800 107.100 88.200 107.200 ;
        RECT 88.600 107.100 89.000 107.200 ;
        RECT 87.800 106.800 89.000 107.100 ;
        RECT 123.800 107.100 124.200 107.200 ;
        RECT 141.400 107.100 141.800 107.200 ;
        RECT 123.800 106.800 141.800 107.100 ;
        RECT 3.800 106.100 4.200 106.200 ;
        RECT 7.800 106.100 8.200 106.200 ;
        RECT 3.800 105.800 8.200 106.100 ;
        RECT 17.400 106.100 17.800 106.200 ;
        RECT 20.600 106.100 21.000 106.200 ;
        RECT 17.400 105.800 21.000 106.100 ;
        RECT 35.000 105.800 35.400 106.200 ;
        RECT 37.400 106.100 37.800 106.200 ;
        RECT 38.200 106.100 38.600 106.200 ;
        RECT 37.400 105.800 38.600 106.100 ;
        RECT 40.600 106.100 41.000 106.200 ;
        RECT 42.200 106.100 42.600 106.200 ;
        RECT 45.400 106.100 45.800 106.200 ;
        RECT 40.600 105.800 45.800 106.100 ;
        RECT 47.000 106.100 47.400 106.200 ;
        RECT 47.800 106.100 48.200 106.200 ;
        RECT 47.000 105.800 48.200 106.100 ;
        RECT 53.400 106.100 53.800 106.200 ;
        RECT 58.200 106.100 58.600 106.200 ;
        RECT 63.000 106.100 63.400 106.200 ;
        RECT 67.800 106.100 68.100 106.800 ;
        RECT 53.400 105.800 60.100 106.100 ;
        RECT 63.000 105.800 68.100 106.100 ;
        RECT 69.400 105.800 69.800 106.200 ;
        RECT 70.200 106.100 70.600 106.200 ;
        RECT 74.200 106.100 74.600 106.200 ;
        RECT 75.800 106.100 76.200 106.200 ;
        RECT 70.200 105.800 76.200 106.100 ;
        RECT 82.200 106.100 82.600 106.200 ;
        RECT 83.000 106.100 83.400 106.200 ;
        RECT 82.200 105.800 83.400 106.100 ;
        RECT 91.800 106.100 92.200 106.200 ;
        RECT 93.400 106.100 93.800 106.200 ;
        RECT 91.800 105.800 93.800 106.100 ;
        RECT 142.200 106.100 142.600 106.200 ;
        RECT 143.000 106.100 143.400 106.200 ;
        RECT 142.200 105.800 143.400 106.100 ;
        RECT 146.200 106.100 146.600 106.200 ;
        RECT 147.000 106.100 147.400 106.200 ;
        RECT 146.200 105.800 147.400 106.100 ;
        RECT 0.600 105.100 1.000 105.200 ;
        RECT 1.400 105.100 1.800 105.200 ;
        RECT 0.600 104.800 1.800 105.100 ;
        RECT 2.200 104.800 2.600 105.200 ;
        RECT 6.200 105.100 6.600 105.200 ;
        RECT 8.600 105.100 9.000 105.200 ;
        RECT 6.200 104.800 9.000 105.100 ;
        RECT 15.000 105.100 15.400 105.200 ;
        RECT 18.200 105.100 18.600 105.200 ;
        RECT 15.000 104.800 18.600 105.100 ;
        RECT 29.400 105.100 29.800 105.200 ;
        RECT 31.800 105.100 32.200 105.200 ;
        RECT 29.400 104.800 32.200 105.100 ;
        RECT 35.000 105.100 35.300 105.800 ;
        RECT 59.800 105.200 60.100 105.800 ;
        RECT 38.200 105.100 38.600 105.200 ;
        RECT 35.000 104.800 38.600 105.100 ;
        RECT 43.000 105.100 43.400 105.200 ;
        RECT 45.400 105.100 45.800 105.200 ;
        RECT 43.000 104.800 45.800 105.100 ;
        RECT 55.000 104.800 55.400 105.200 ;
        RECT 59.800 104.800 60.200 105.200 ;
        RECT 63.000 105.100 63.400 105.200 ;
        RECT 63.800 105.100 64.200 105.200 ;
        RECT 63.000 104.800 64.200 105.100 ;
        RECT 64.600 105.100 65.000 105.200 ;
        RECT 65.400 105.100 65.800 105.200 ;
        RECT 64.600 104.800 65.800 105.100 ;
        RECT 67.000 105.100 67.400 105.200 ;
        RECT 69.400 105.100 69.700 105.800 ;
        RECT 67.000 104.800 69.700 105.100 ;
        RECT 72.600 105.100 73.000 105.200 ;
        RECT 75.000 105.100 75.400 105.200 ;
        RECT 83.000 105.100 83.400 105.200 ;
        RECT 72.600 104.800 83.400 105.100 ;
        RECT 115.800 105.100 116.200 105.200 ;
        RECT 119.800 105.100 120.200 105.200 ;
        RECT 115.800 104.800 120.200 105.100 ;
        RECT 139.800 105.100 140.200 105.200 ;
        RECT 142.200 105.100 142.600 105.200 ;
        RECT 139.800 104.800 142.600 105.100 ;
        RECT 2.200 104.100 2.500 104.800 ;
        RECT 19.800 104.100 20.200 104.200 ;
        RECT 2.200 103.800 20.200 104.100 ;
        RECT 21.400 104.100 21.800 104.200 ;
        RECT 23.000 104.100 23.400 104.200 ;
        RECT 21.400 103.800 23.400 104.100 ;
        RECT 26.200 104.100 26.600 104.200 ;
        RECT 31.000 104.100 31.400 104.200 ;
        RECT 31.800 104.100 32.200 104.200 ;
        RECT 26.200 103.800 32.200 104.100 ;
        RECT 32.600 104.100 33.000 104.200 ;
        RECT 40.600 104.100 41.000 104.200 ;
        RECT 32.600 103.800 41.000 104.100 ;
        RECT 42.200 104.100 42.600 104.200 ;
        RECT 47.800 104.100 48.200 104.200 ;
        RECT 55.000 104.100 55.300 104.800 ;
        RECT 42.200 103.800 55.300 104.100 ;
        RECT 55.800 104.100 56.200 104.200 ;
        RECT 59.000 104.100 59.400 104.200 ;
        RECT 62.200 104.100 62.600 104.200 ;
        RECT 55.800 103.800 62.600 104.100 ;
        RECT 81.400 104.100 81.800 104.200 ;
        RECT 85.400 104.100 85.800 104.200 ;
        RECT 91.000 104.100 91.400 104.200 ;
        RECT 81.400 103.800 91.400 104.100 ;
        RECT 115.000 104.100 115.400 104.200 ;
        RECT 124.600 104.100 125.000 104.200 ;
        RECT 115.000 103.800 125.000 104.100 ;
        RECT 2.200 102.800 2.600 103.200 ;
        RECT 22.200 103.100 22.600 103.200 ;
        RECT 24.600 103.100 25.000 103.200 ;
        RECT 22.200 102.800 25.000 103.100 ;
        RECT 27.800 103.100 28.200 103.200 ;
        RECT 30.200 103.100 30.600 103.200 ;
        RECT 33.400 103.100 33.800 103.200 ;
        RECT 46.200 103.100 46.600 103.200 ;
        RECT 27.800 102.800 46.600 103.100 ;
        RECT 51.800 103.100 52.200 103.200 ;
        RECT 53.400 103.100 53.800 103.200 ;
        RECT 69.400 103.100 69.800 103.200 ;
        RECT 51.800 102.800 69.800 103.100 ;
        RECT 87.800 103.100 88.200 103.200 ;
        RECT 122.200 103.100 122.600 103.200 ;
        RECT 87.800 102.800 122.600 103.100 ;
        RECT 2.200 102.200 2.500 102.800 ;
        RECT 2.200 101.800 2.600 102.200 ;
        RECT 55.800 102.100 56.200 102.200 ;
        RECT 65.400 102.100 65.800 102.200 ;
        RECT 55.800 101.800 65.800 102.100 ;
        RECT 79.800 102.100 80.200 102.200 ;
        RECT 83.800 102.100 84.200 102.200 ;
        RECT 87.800 102.100 88.200 102.200 ;
        RECT 79.800 101.800 88.200 102.100 ;
        RECT 119.800 102.100 120.200 102.200 ;
        RECT 121.400 102.100 121.800 102.200 ;
        RECT 119.800 101.800 121.800 102.100 ;
        RECT 51.000 101.100 51.400 101.200 ;
        RECT 59.000 101.100 59.400 101.200 ;
        RECT 51.000 100.800 59.400 101.100 ;
        RECT 99.000 101.100 99.400 101.200 ;
        RECT 106.200 101.100 106.600 101.200 ;
        RECT 99.000 100.800 106.600 101.100 ;
        RECT 7.800 99.100 8.200 99.200 ;
        RECT 10.200 99.100 10.600 99.200 ;
        RECT 7.800 98.800 10.600 99.100 ;
        RECT 45.400 99.100 45.800 99.200 ;
        RECT 51.800 99.100 52.200 99.200 ;
        RECT 45.400 98.800 52.200 99.100 ;
        RECT 82.200 99.100 82.600 99.200 ;
        RECT 86.200 99.100 86.600 99.200 ;
        RECT 82.200 98.800 86.600 99.100 ;
        RECT 87.000 99.100 87.400 99.200 ;
        RECT 97.400 99.100 97.800 99.200 ;
        RECT 87.000 98.800 97.800 99.100 ;
        RECT 109.400 99.100 109.800 99.200 ;
        RECT 119.800 99.100 120.200 99.200 ;
        RECT 109.400 98.800 120.200 99.100 ;
        RECT 26.200 98.100 26.600 98.200 ;
        RECT 28.600 98.100 29.000 98.200 ;
        RECT 31.800 98.100 32.200 98.200 ;
        RECT 38.200 98.100 38.600 98.200 ;
        RECT 26.200 97.800 38.600 98.100 ;
        RECT 40.600 97.800 41.000 98.200 ;
        RECT 47.000 98.100 47.400 98.200 ;
        RECT 51.800 98.100 52.200 98.200 ;
        RECT 47.000 97.800 52.200 98.100 ;
        RECT 77.400 98.100 77.800 98.200 ;
        RECT 89.400 98.100 89.800 98.200 ;
        RECT 77.400 97.800 89.800 98.100 ;
        RECT 96.600 98.100 97.000 98.200 ;
        RECT 105.400 98.100 105.800 98.200 ;
        RECT 96.600 97.800 105.800 98.100 ;
        RECT 2.200 97.100 2.600 97.200 ;
        RECT 5.400 97.100 5.800 97.200 ;
        RECT 6.200 97.100 6.600 97.200 ;
        RECT 2.200 96.800 6.600 97.100 ;
        RECT 8.600 97.100 9.000 97.200 ;
        RECT 16.600 97.100 17.000 97.200 ;
        RECT 19.000 97.100 19.400 97.200 ;
        RECT 8.600 96.800 19.400 97.100 ;
        RECT 34.200 97.100 34.600 97.200 ;
        RECT 39.800 97.100 40.200 97.200 ;
        RECT 40.600 97.100 40.900 97.800 ;
        RECT 43.000 97.100 43.400 97.200 ;
        RECT 34.200 96.800 43.400 97.100 ;
        RECT 46.200 97.100 46.600 97.200 ;
        RECT 51.000 97.100 51.400 97.200 ;
        RECT 54.200 97.100 54.600 97.200 ;
        RECT 46.200 96.800 54.600 97.100 ;
        RECT 65.400 97.100 65.800 97.200 ;
        RECT 71.000 97.100 71.400 97.200 ;
        RECT 79.000 97.100 79.400 97.200 ;
        RECT 65.400 96.800 79.400 97.100 ;
        RECT 87.000 97.100 87.400 97.200 ;
        RECT 95.000 97.100 95.400 97.200 ;
        RECT 87.000 96.800 95.400 97.100 ;
        RECT 99.000 96.800 99.400 97.200 ;
        RECT 9.400 96.100 9.800 96.200 ;
        RECT 15.800 96.100 16.200 96.200 ;
        RECT 20.600 96.100 21.000 96.200 ;
        RECT 9.400 95.800 21.000 96.100 ;
        RECT 23.000 96.100 23.400 96.200 ;
        RECT 23.800 96.100 24.200 96.200 ;
        RECT 23.000 95.800 24.200 96.100 ;
        RECT 37.400 96.100 37.800 96.200 ;
        RECT 54.200 96.100 54.600 96.200 ;
        RECT 37.400 95.800 54.600 96.100 ;
        RECT 67.800 96.100 68.200 96.200 ;
        RECT 69.400 96.100 69.800 96.200 ;
        RECT 67.800 95.800 69.800 96.100 ;
        RECT 74.200 96.100 74.600 96.200 ;
        RECT 76.600 96.100 77.000 96.200 ;
        RECT 87.000 96.100 87.400 96.200 ;
        RECT 74.200 95.800 87.400 96.100 ;
        RECT 96.600 96.100 97.000 96.200 ;
        RECT 99.000 96.100 99.300 96.800 ;
        RECT 139.900 96.100 140.300 96.200 ;
        RECT 96.600 95.800 99.300 96.100 ;
        RECT 139.800 95.800 140.300 96.100 ;
        RECT 4.600 95.100 5.000 95.200 ;
        RECT 6.200 95.100 6.600 95.200 ;
        RECT 4.600 94.800 6.600 95.100 ;
        RECT 29.400 95.100 29.800 95.200 ;
        RECT 31.800 95.100 32.200 95.200 ;
        RECT 29.400 94.800 32.200 95.100 ;
        RECT 35.000 94.800 35.400 95.200 ;
        RECT 35.800 95.100 36.200 95.200 ;
        RECT 39.000 95.100 39.400 95.200 ;
        RECT 52.600 95.100 53.000 95.200 ;
        RECT 35.800 94.800 53.000 95.100 ;
        RECT 62.200 95.100 62.600 95.200 ;
        RECT 71.800 95.100 72.200 95.200 ;
        RECT 62.200 94.800 72.200 95.100 ;
        RECT 75.800 95.100 76.200 95.200 ;
        RECT 76.600 95.100 77.000 95.200 ;
        RECT 75.800 94.800 77.000 95.100 ;
        RECT 77.400 95.100 77.800 95.200 ;
        RECT 79.000 95.100 79.400 95.200 ;
        RECT 77.400 94.800 79.400 95.100 ;
        RECT 80.600 95.100 81.000 95.200 ;
        RECT 81.400 95.100 81.800 95.200 ;
        RECT 91.800 95.100 92.200 95.200 ;
        RECT 80.600 94.800 81.800 95.100 ;
        RECT 82.200 94.800 92.200 95.100 ;
        RECT 99.000 95.100 99.400 95.200 ;
        RECT 107.000 95.100 107.400 95.200 ;
        RECT 99.000 94.800 107.400 95.100 ;
        RECT 118.200 94.800 118.600 95.200 ;
        RECT 139.800 95.100 140.100 95.800 ;
        RECT 143.800 95.100 144.200 95.200 ;
        RECT 147.000 95.100 147.400 95.200 ;
        RECT 139.800 94.800 147.400 95.100 ;
        RECT 148.600 94.800 149.000 95.200 ;
        RECT 0.600 94.100 1.000 94.200 ;
        RECT 3.000 94.100 3.400 94.200 ;
        RECT 22.200 94.100 22.600 94.200 ;
        RECT 0.600 93.800 3.400 94.100 ;
        RECT 12.600 93.800 22.600 94.100 ;
        RECT 24.600 94.100 25.000 94.200 ;
        RECT 35.000 94.100 35.300 94.800 ;
        RECT 24.600 93.800 35.300 94.100 ;
        RECT 36.600 94.100 37.000 94.200 ;
        RECT 37.400 94.100 37.800 94.200 ;
        RECT 36.600 93.800 37.800 94.100 ;
        RECT 39.000 94.100 39.400 94.200 ;
        RECT 40.600 94.100 41.000 94.200 ;
        RECT 39.000 93.800 41.000 94.100 ;
        RECT 42.200 94.100 42.600 94.200 ;
        RECT 53.400 94.100 53.800 94.200 ;
        RECT 55.000 94.100 55.400 94.200 ;
        RECT 42.200 93.800 55.400 94.100 ;
        RECT 59.800 94.100 60.200 94.200 ;
        RECT 64.600 94.100 65.000 94.200 ;
        RECT 67.000 94.100 67.400 94.200 ;
        RECT 59.800 93.800 64.100 94.100 ;
        RECT 64.600 93.800 67.400 94.100 ;
        RECT 72.600 94.100 73.000 94.200 ;
        RECT 73.400 94.100 73.800 94.200 ;
        RECT 72.600 93.800 73.800 94.100 ;
        RECT 77.400 94.100 77.800 94.200 ;
        RECT 78.200 94.100 78.600 94.200 ;
        RECT 82.200 94.100 82.500 94.800 ;
        RECT 118.200 94.200 118.500 94.800 ;
        RECT 148.600 94.200 148.900 94.800 ;
        RECT 77.400 93.800 82.500 94.100 ;
        RECT 92.600 94.100 93.000 94.200 ;
        RECT 96.600 94.100 97.000 94.200 ;
        RECT 92.600 93.800 97.000 94.100 ;
        RECT 103.000 94.100 103.400 94.200 ;
        RECT 103.800 94.100 104.200 94.200 ;
        RECT 103.000 93.800 104.200 94.100 ;
        RECT 105.400 94.100 105.800 94.200 ;
        RECT 110.200 94.100 110.600 94.200 ;
        RECT 105.400 93.800 110.600 94.100 ;
        RECT 114.200 93.800 114.600 94.200 ;
        RECT 118.200 93.800 118.600 94.200 ;
        RECT 119.000 94.100 119.400 94.200 ;
        RECT 119.800 94.100 120.200 94.200 ;
        RECT 119.000 93.800 120.200 94.100 ;
        RECT 122.200 94.100 122.600 94.200 ;
        RECT 139.800 94.100 140.200 94.200 ;
        RECT 122.200 93.800 140.200 94.100 ;
        RECT 148.600 93.800 149.000 94.200 ;
        RECT 12.600 93.200 12.900 93.800 ;
        RECT 63.800 93.200 64.100 93.800 ;
        RECT 114.200 93.200 114.500 93.800 ;
        RECT 2.200 93.100 2.600 93.200 ;
        RECT 8.600 93.100 9.000 93.200 ;
        RECT 11.800 93.100 12.200 93.200 ;
        RECT 2.200 92.800 12.200 93.100 ;
        RECT 12.600 92.800 13.000 93.200 ;
        RECT 25.400 92.800 25.800 93.200 ;
        RECT 27.000 93.100 27.400 93.200 ;
        RECT 30.200 93.100 30.600 93.200 ;
        RECT 50.200 93.100 50.600 93.200 ;
        RECT 27.000 92.800 50.600 93.100 ;
        RECT 63.800 92.800 64.200 93.200 ;
        RECT 72.600 93.100 73.000 93.200 ;
        RECT 75.000 93.100 75.400 93.200 ;
        RECT 83.000 93.100 83.400 93.200 ;
        RECT 72.600 92.800 83.400 93.100 ;
        RECT 93.400 93.100 93.800 93.200 ;
        RECT 94.200 93.100 94.600 93.200 ;
        RECT 99.000 93.100 99.400 93.200 ;
        RECT 93.400 92.800 99.400 93.100 ;
        RECT 103.000 93.100 103.400 93.200 ;
        RECT 103.800 93.100 104.200 93.200 ;
        RECT 103.000 92.800 104.200 93.100 ;
        RECT 114.200 92.800 114.600 93.200 ;
        RECT 122.200 93.100 122.600 93.200 ;
        RECT 145.400 93.100 145.800 93.200 ;
        RECT 122.200 92.800 145.800 93.100 ;
        RECT 3.800 92.100 4.200 92.200 ;
        RECT 4.600 92.100 5.000 92.200 ;
        RECT 3.800 91.800 5.000 92.100 ;
        RECT 10.200 92.100 10.600 92.200 ;
        RECT 25.400 92.100 25.700 92.800 ;
        RECT 10.200 91.800 25.700 92.100 ;
        RECT 33.400 92.100 33.800 92.200 ;
        RECT 43.800 92.100 44.200 92.200 ;
        RECT 45.400 92.100 45.800 92.200 ;
        RECT 33.400 91.800 45.800 92.100 ;
        RECT 52.600 92.100 53.000 92.200 ;
        RECT 55.000 92.100 55.400 92.200 ;
        RECT 52.600 91.800 55.400 92.100 ;
        RECT 60.600 92.100 61.000 92.200 ;
        RECT 64.600 92.100 65.000 92.200 ;
        RECT 60.600 91.800 65.000 92.100 ;
        RECT 71.000 92.100 71.400 92.200 ;
        RECT 76.600 92.100 77.000 92.200 ;
        RECT 71.000 91.800 77.000 92.100 ;
        RECT 80.600 92.100 81.000 92.200 ;
        RECT 83.800 92.100 84.200 92.200 ;
        RECT 80.600 91.800 84.200 92.100 ;
        RECT 84.600 92.100 85.000 92.200 ;
        RECT 91.000 92.100 91.400 92.200 ;
        RECT 84.600 91.800 91.400 92.100 ;
        RECT 98.200 92.100 98.600 92.200 ;
        RECT 109.400 92.100 109.800 92.200 ;
        RECT 98.200 91.800 109.800 92.100 ;
        RECT 115.800 92.100 116.200 92.200 ;
        RECT 124.600 92.100 125.000 92.200 ;
        RECT 115.800 91.800 125.000 92.100 ;
        RECT 14.200 90.800 14.600 91.200 ;
        RECT 15.800 91.100 16.200 91.200 ;
        RECT 25.400 91.100 25.800 91.200 ;
        RECT 15.800 90.800 25.800 91.100 ;
        RECT 63.800 91.100 64.200 91.200 ;
        RECT 65.400 91.100 65.800 91.200 ;
        RECT 63.800 90.800 65.800 91.100 ;
        RECT 69.400 91.100 69.800 91.200 ;
        RECT 71.800 91.100 72.200 91.200 ;
        RECT 69.400 90.800 72.200 91.100 ;
        RECT 14.200 90.200 14.500 90.800 ;
        RECT 14.200 89.800 14.600 90.200 ;
        RECT 81.400 90.100 81.800 90.200 ;
        RECT 88.600 90.100 89.000 90.200 ;
        RECT 109.400 90.100 109.800 90.200 ;
        RECT 113.400 90.100 113.800 90.200 ;
        RECT 128.600 90.100 129.000 90.200 ;
        RECT 81.400 89.800 94.500 90.100 ;
        RECT 109.400 89.800 129.000 90.100 ;
        RECT 1.400 89.100 1.800 89.200 ;
        RECT 7.000 89.100 7.400 89.200 ;
        RECT 1.400 88.800 7.400 89.100 ;
        RECT 15.800 89.100 16.200 89.200 ;
        RECT 21.400 89.100 21.800 89.200 ;
        RECT 15.800 88.800 21.800 89.100 ;
        RECT 37.400 89.100 37.800 89.200 ;
        RECT 41.400 89.100 41.800 89.200 ;
        RECT 37.400 88.800 41.800 89.100 ;
        RECT 44.600 89.100 45.000 89.200 ;
        RECT 54.200 89.100 54.600 89.200 ;
        RECT 44.600 88.800 54.600 89.100 ;
        RECT 63.000 89.100 63.400 89.200 ;
        RECT 74.200 89.100 74.600 89.200 ;
        RECT 63.000 88.800 74.600 89.100 ;
        RECT 87.000 88.800 87.400 89.200 ;
        RECT 87.800 89.100 88.200 89.200 ;
        RECT 93.400 89.100 93.800 89.200 ;
        RECT 87.800 88.800 93.800 89.100 ;
        RECT 94.200 89.100 94.500 89.800 ;
        RECT 94.200 88.800 106.500 89.100 ;
        RECT 7.800 88.100 8.200 88.200 ;
        RECT 10.200 88.100 10.600 88.200 ;
        RECT 7.800 87.800 10.600 88.100 ;
        RECT 30.200 88.100 30.600 88.200 ;
        RECT 40.600 88.100 41.000 88.200 ;
        RECT 56.600 88.100 57.000 88.200 ;
        RECT 30.200 87.800 57.000 88.100 ;
        RECT 57.400 87.800 57.800 88.200 ;
        RECT 59.000 88.100 59.400 88.200 ;
        RECT 61.400 88.100 61.800 88.200 ;
        RECT 63.800 88.100 64.200 88.200 ;
        RECT 59.000 87.800 64.200 88.100 ;
        RECT 87.000 88.100 87.300 88.800 ;
        RECT 106.200 88.200 106.500 88.800 ;
        RECT 119.800 88.800 120.200 89.200 ;
        RECT 130.200 89.100 130.600 89.200 ;
        RECT 140.600 89.100 141.000 89.200 ;
        RECT 130.200 88.800 141.000 89.100 ;
        RECT 94.200 88.100 94.600 88.200 ;
        RECT 87.000 87.800 94.600 88.100 ;
        RECT 106.200 87.800 106.600 88.200 ;
        RECT 118.200 88.100 118.600 88.200 ;
        RECT 119.800 88.100 120.100 88.800 ;
        RECT 118.200 87.800 120.100 88.100 ;
        RECT 123.800 88.100 124.200 88.200 ;
        RECT 124.600 88.100 125.000 88.200 ;
        RECT 126.200 88.100 126.600 88.200 ;
        RECT 131.000 88.100 131.400 88.200 ;
        RECT 123.800 87.800 131.400 88.100 ;
        RECT 143.800 88.100 144.200 88.200 ;
        RECT 144.600 88.100 145.000 88.200 ;
        RECT 143.800 87.800 145.000 88.100 ;
        RECT 7.000 87.100 7.400 87.200 ;
        RECT 7.800 87.100 8.200 87.200 ;
        RECT 7.000 86.800 8.200 87.100 ;
        RECT 8.600 87.100 9.000 87.200 ;
        RECT 12.600 87.100 13.000 87.200 ;
        RECT 17.400 87.100 17.800 87.200 ;
        RECT 8.600 86.800 17.800 87.100 ;
        RECT 25.400 87.100 25.800 87.200 ;
        RECT 27.000 87.100 27.400 87.200 ;
        RECT 25.400 86.800 27.400 87.100 ;
        RECT 34.200 87.100 34.600 87.200 ;
        RECT 38.200 87.100 38.600 87.200 ;
        RECT 34.200 86.800 38.600 87.100 ;
        RECT 39.800 87.100 40.200 87.200 ;
        RECT 40.600 87.100 41.000 87.200 ;
        RECT 43.000 87.100 43.400 87.200 ;
        RECT 39.800 86.800 43.400 87.100 ;
        RECT 48.600 87.100 49.000 87.200 ;
        RECT 53.400 87.100 53.800 87.200 ;
        RECT 57.400 87.100 57.700 87.800 ;
        RECT 48.600 86.800 57.700 87.100 ;
        RECT 89.400 86.800 89.800 87.200 ;
        RECT 91.000 87.100 91.400 87.200 ;
        RECT 106.200 87.100 106.600 87.200 ;
        RECT 91.000 86.800 106.600 87.100 ;
        RECT 107.800 87.100 108.200 87.200 ;
        RECT 109.400 87.100 109.800 87.200 ;
        RECT 107.800 86.800 109.800 87.100 ;
        RECT 111.000 86.800 111.400 87.200 ;
        RECT 111.800 87.100 112.200 87.200 ;
        RECT 115.800 87.100 116.200 87.200 ;
        RECT 111.800 86.800 116.200 87.100 ;
        RECT 122.200 87.100 122.600 87.200 ;
        RECT 123.800 87.100 124.200 87.200 ;
        RECT 122.200 86.800 124.200 87.100 ;
        RECT 125.400 87.100 125.800 87.200 ;
        RECT 130.200 87.100 130.600 87.200 ;
        RECT 131.800 87.100 132.200 87.200 ;
        RECT 125.400 86.800 128.100 87.100 ;
        RECT 130.200 86.800 132.200 87.100 ;
        RECT 3.000 86.100 3.400 86.200 ;
        RECT 4.600 86.100 5.000 86.200 ;
        RECT 9.400 86.100 9.800 86.200 ;
        RECT 3.000 85.800 9.800 86.100 ;
        RECT 14.200 86.100 14.600 86.200 ;
        RECT 18.200 86.100 18.600 86.200 ;
        RECT 14.200 85.800 18.600 86.100 ;
        RECT 27.800 86.100 28.200 86.200 ;
        RECT 32.600 86.100 33.000 86.200 ;
        RECT 27.800 85.800 33.000 86.100 ;
        RECT 34.200 85.800 34.600 86.200 ;
        RECT 39.000 86.100 39.400 86.200 ;
        RECT 35.800 85.800 39.400 86.100 ;
        RECT 63.800 85.800 64.200 86.200 ;
        RECT 75.800 86.100 76.200 86.200 ;
        RECT 81.400 86.100 81.800 86.200 ;
        RECT 89.400 86.100 89.700 86.800 ;
        RECT 75.800 85.800 89.700 86.100 ;
        RECT 103.800 85.800 104.200 86.200 ;
        RECT 111.000 86.100 111.300 86.800 ;
        RECT 127.800 86.200 128.100 86.800 ;
        RECT 117.400 86.100 117.800 86.200 ;
        RECT 119.000 86.100 119.400 86.200 ;
        RECT 123.000 86.100 123.400 86.200 ;
        RECT 126.200 86.100 126.600 86.200 ;
        RECT 111.000 85.800 126.600 86.100 ;
        RECT 127.800 85.800 128.200 86.200 ;
        RECT 139.000 86.100 139.400 86.200 ;
        RECT 135.800 85.800 139.400 86.100 ;
        RECT 0.600 85.100 1.000 85.200 ;
        RECT 15.000 85.100 15.400 85.200 ;
        RECT 0.600 84.800 15.400 85.100 ;
        RECT 19.800 85.100 20.200 85.200 ;
        RECT 25.400 85.100 25.800 85.200 ;
        RECT 28.600 85.100 29.000 85.200 ;
        RECT 19.800 84.800 29.000 85.100 ;
        RECT 29.400 85.100 29.800 85.200 ;
        RECT 31.800 85.100 32.200 85.200 ;
        RECT 34.200 85.100 34.500 85.800 ;
        RECT 29.400 84.800 34.500 85.100 ;
        RECT 35.800 85.200 36.100 85.800 ;
        RECT 39.000 85.200 39.300 85.800 ;
        RECT 35.800 84.800 36.200 85.200 ;
        RECT 39.000 84.800 39.400 85.200 ;
        RECT 41.400 85.100 41.800 85.200 ;
        RECT 43.800 85.100 44.200 85.200 ;
        RECT 44.600 85.100 45.000 85.200 ;
        RECT 41.400 84.800 45.000 85.100 ;
        RECT 45.400 85.100 45.800 85.200 ;
        RECT 47.800 85.100 48.200 85.200 ;
        RECT 52.600 85.100 53.000 85.200 ;
        RECT 45.400 84.800 53.000 85.100 ;
        RECT 53.400 84.800 53.800 85.200 ;
        RECT 56.600 85.100 57.000 85.200 ;
        RECT 63.800 85.100 64.100 85.800 ;
        RECT 103.800 85.200 104.100 85.800 ;
        RECT 135.800 85.200 136.100 85.800 ;
        RECT 56.600 84.800 64.100 85.100 ;
        RECT 66.200 85.100 66.600 85.200 ;
        RECT 87.000 85.100 87.400 85.200 ;
        RECT 66.200 84.800 87.400 85.100 ;
        RECT 103.800 84.800 104.200 85.200 ;
        RECT 135.800 84.800 136.200 85.200 ;
        RECT 137.400 85.100 137.800 85.200 ;
        RECT 137.400 84.800 146.500 85.100 ;
        RECT 8.600 84.100 9.000 84.200 ;
        RECT 19.000 84.100 19.400 84.200 ;
        RECT 35.800 84.100 36.200 84.200 ;
        RECT 39.800 84.100 40.200 84.200 ;
        RECT 8.600 83.800 32.900 84.100 ;
        RECT 35.800 83.800 40.200 84.100 ;
        RECT 51.800 84.100 52.200 84.200 ;
        RECT 53.400 84.100 53.700 84.800 ;
        RECT 146.200 84.200 146.500 84.800 ;
        RECT 51.800 83.800 53.700 84.100 ;
        RECT 59.800 84.100 60.200 84.200 ;
        RECT 64.600 84.100 65.000 84.200 ;
        RECT 59.800 83.800 65.000 84.100 ;
        RECT 67.000 84.100 67.400 84.200 ;
        RECT 68.600 84.100 69.000 84.200 ;
        RECT 67.000 83.800 69.000 84.100 ;
        RECT 114.200 84.100 114.600 84.200 ;
        RECT 135.800 84.100 136.200 84.200 ;
        RECT 138.200 84.100 138.600 84.200 ;
        RECT 114.200 83.800 138.600 84.100 ;
        RECT 146.200 84.100 146.600 84.200 ;
        RECT 150.200 84.100 150.600 84.200 ;
        RECT 146.200 83.800 150.600 84.100 ;
        RECT 32.600 83.200 32.900 83.800 ;
        RECT 32.600 82.800 33.000 83.200 ;
        RECT 87.000 83.100 87.400 83.200 ;
        RECT 91.000 83.100 91.400 83.200 ;
        RECT 93.400 83.100 93.800 83.200 ;
        RECT 87.000 82.800 93.800 83.100 ;
        RECT 128.600 83.100 129.000 83.200 ;
        RECT 139.000 83.100 139.400 83.200 ;
        RECT 128.600 82.800 139.400 83.100 ;
        RECT 9.400 82.100 9.800 82.200 ;
        RECT 12.600 82.100 13.000 82.200 ;
        RECT 16.600 82.100 17.000 82.200 ;
        RECT 17.400 82.100 17.800 82.200 ;
        RECT 9.400 81.800 17.800 82.100 ;
        RECT 81.400 82.100 81.800 82.200 ;
        RECT 83.800 82.100 84.200 82.200 ;
        RECT 81.400 81.800 84.200 82.100 ;
        RECT 87.800 82.100 88.200 82.200 ;
        RECT 95.800 82.100 96.200 82.200 ;
        RECT 87.800 81.800 96.200 82.100 ;
        RECT 96.600 82.100 97.000 82.200 ;
        RECT 108.600 82.100 109.000 82.200 ;
        RECT 96.600 81.800 109.000 82.100 ;
        RECT 123.800 82.100 124.200 82.200 ;
        RECT 148.600 82.100 149.000 82.200 ;
        RECT 123.800 81.800 149.000 82.100 ;
        RECT 17.400 80.800 17.800 81.200 ;
        RECT 53.400 81.100 53.800 81.200 ;
        RECT 55.000 81.100 55.400 81.200 ;
        RECT 53.400 80.800 55.400 81.100 ;
        RECT 73.400 81.100 73.800 81.200 ;
        RECT 75.800 81.100 76.200 81.200 ;
        RECT 73.400 80.800 76.200 81.100 ;
        RECT 77.400 80.800 77.800 81.200 ;
        RECT 87.800 81.100 88.200 81.200 ;
        RECT 112.600 81.100 113.000 81.200 ;
        RECT 87.800 80.800 113.000 81.100 ;
        RECT 17.400 80.200 17.700 80.800 ;
        RECT 77.400 80.200 77.700 80.800 ;
        RECT 17.400 79.800 17.800 80.200 ;
        RECT 51.000 80.100 51.400 80.200 ;
        RECT 55.800 80.100 56.200 80.200 ;
        RECT 51.000 79.800 56.200 80.100 ;
        RECT 63.000 80.100 63.400 80.200 ;
        RECT 72.600 80.100 73.000 80.200 ;
        RECT 75.000 80.100 75.400 80.200 ;
        RECT 63.000 79.800 75.400 80.100 ;
        RECT 77.400 79.800 77.800 80.200 ;
        RECT 81.400 80.100 81.800 80.200 ;
        RECT 107.800 80.100 108.200 80.200 ;
        RECT 110.200 80.100 110.600 80.200 ;
        RECT 81.400 79.800 110.600 80.100 ;
        RECT 119.000 80.100 119.400 80.200 ;
        RECT 135.800 80.100 136.200 80.200 ;
        RECT 119.000 79.800 136.200 80.100 ;
        RECT 3.800 79.100 4.200 79.200 ;
        RECT 5.400 79.100 5.800 79.200 ;
        RECT 3.800 78.800 5.800 79.100 ;
        RECT 7.800 79.100 8.200 79.200 ;
        RECT 14.200 79.100 14.600 79.200 ;
        RECT 7.800 78.800 14.600 79.100 ;
        RECT 27.000 79.100 27.400 79.200 ;
        RECT 59.800 79.100 60.200 79.200 ;
        RECT 27.000 78.800 60.200 79.100 ;
        RECT 71.800 79.100 72.200 79.200 ;
        RECT 73.400 79.100 73.800 79.200 ;
        RECT 102.200 79.100 102.600 79.200 ;
        RECT 71.800 78.800 73.800 79.100 ;
        RECT 82.200 78.800 102.600 79.100 ;
        RECT 107.000 79.100 107.400 79.200 ;
        RECT 122.200 79.100 122.600 79.200 ;
        RECT 127.000 79.100 127.400 79.200 ;
        RECT 131.000 79.100 131.400 79.200 ;
        RECT 131.800 79.100 132.200 79.200 ;
        RECT 107.000 78.800 132.200 79.100 ;
        RECT 82.200 78.200 82.500 78.800 ;
        RECT 45.400 78.100 45.800 78.200 ;
        RECT 49.400 78.100 49.800 78.200 ;
        RECT 45.400 77.800 52.900 78.100 ;
        RECT 52.600 77.200 52.900 77.800 ;
        RECT 55.800 77.800 56.200 78.200 ;
        RECT 61.400 78.100 61.800 78.200 ;
        RECT 74.200 78.100 74.600 78.200 ;
        RECT 80.600 78.100 81.000 78.200 ;
        RECT 61.400 77.800 81.000 78.100 ;
        RECT 82.200 77.800 82.600 78.200 ;
        RECT 89.400 78.100 89.800 78.200 ;
        RECT 94.200 78.100 94.600 78.200 ;
        RECT 136.600 78.100 137.000 78.200 ;
        RECT 89.400 77.800 94.600 78.100 ;
        RECT 128.600 77.800 137.000 78.100 ;
        RECT 137.400 77.800 137.800 78.200 ;
        RECT 19.800 76.800 20.200 77.200 ;
        RECT 33.400 76.800 33.800 77.200 ;
        RECT 43.000 77.100 43.400 77.200 ;
        RECT 50.200 77.100 50.600 77.200 ;
        RECT 43.000 76.800 50.600 77.100 ;
        RECT 52.600 76.800 53.000 77.200 ;
        RECT 55.800 77.100 56.100 77.800 ;
        RECT 128.600 77.200 128.900 77.800 ;
        RECT 58.200 77.100 58.600 77.200 ;
        RECT 55.800 76.800 58.600 77.100 ;
        RECT 68.600 77.100 69.000 77.200 ;
        RECT 75.800 77.100 76.200 77.200 ;
        RECT 87.800 77.100 88.200 77.200 ;
        RECT 68.600 76.800 88.200 77.100 ;
        RECT 88.600 77.100 89.000 77.200 ;
        RECT 91.800 77.100 92.200 77.200 ;
        RECT 92.600 77.100 93.000 77.200 ;
        RECT 88.600 76.800 93.000 77.100 ;
        RECT 95.800 77.100 96.200 77.200 ;
        RECT 107.800 77.100 108.200 77.200 ;
        RECT 120.600 77.100 121.000 77.200 ;
        RECT 95.800 76.800 121.000 77.100 ;
        RECT 121.400 76.800 121.800 77.200 ;
        RECT 128.600 76.800 129.000 77.200 ;
        RECT 132.600 76.800 133.000 77.200 ;
        RECT 134.200 77.100 134.600 77.200 ;
        RECT 137.400 77.100 137.700 77.800 ;
        RECT 134.200 76.800 137.700 77.100 ;
        RECT 3.800 76.100 4.200 76.200 ;
        RECT 6.200 76.100 6.600 76.200 ;
        RECT 3.800 75.800 6.600 76.100 ;
        RECT 10.200 76.100 10.600 76.200 ;
        RECT 12.600 76.100 13.000 76.200 ;
        RECT 10.200 75.800 13.000 76.100 ;
        RECT 17.400 76.100 17.800 76.200 ;
        RECT 19.800 76.100 20.100 76.800 ;
        RECT 17.400 75.800 20.100 76.100 ;
        RECT 25.400 76.100 25.800 76.200 ;
        RECT 27.000 76.100 27.400 76.200 ;
        RECT 33.400 76.100 33.700 76.800 ;
        RECT 25.400 75.800 27.400 76.100 ;
        RECT 27.800 75.800 33.700 76.100 ;
        RECT 84.600 76.100 85.000 76.200 ;
        RECT 85.400 76.100 85.800 76.200 ;
        RECT 94.200 76.100 94.600 76.200 ;
        RECT 84.600 75.800 94.600 76.100 ;
        RECT 95.000 76.100 95.400 76.200 ;
        RECT 97.400 76.100 97.800 76.200 ;
        RECT 98.200 76.100 98.600 76.200 ;
        RECT 95.000 75.800 98.600 76.100 ;
        RECT 99.000 75.800 99.400 76.200 ;
        RECT 114.200 76.100 114.600 76.200 ;
        RECT 121.400 76.100 121.700 76.800 ;
        RECT 129.400 76.100 129.800 76.200 ;
        RECT 114.200 75.800 129.800 76.100 ;
        RECT 130.200 76.100 130.600 76.200 ;
        RECT 131.800 76.100 132.200 76.200 ;
        RECT 130.200 75.800 132.200 76.100 ;
        RECT 132.600 76.100 132.900 76.800 ;
        RECT 136.600 76.100 137.000 76.200 ;
        RECT 137.400 76.100 137.800 76.200 ;
        RECT 132.600 75.800 137.800 76.100 ;
        RECT 139.000 75.800 139.400 76.200 ;
        RECT 145.400 75.800 145.800 76.200 ;
        RECT 6.200 75.100 6.600 75.200 ;
        RECT 7.000 75.100 7.400 75.200 ;
        RECT 9.400 75.100 9.800 75.200 ;
        RECT 6.200 74.800 9.800 75.100 ;
        RECT 20.600 75.100 21.000 75.200 ;
        RECT 23.000 75.100 23.400 75.200 ;
        RECT 20.600 74.800 23.400 75.100 ;
        RECT 27.000 75.100 27.400 75.200 ;
        RECT 27.800 75.100 28.100 75.800 ;
        RECT 99.000 75.200 99.300 75.800 ;
        RECT 139.000 75.200 139.300 75.800 ;
        RECT 27.000 74.800 28.100 75.100 ;
        RECT 50.200 75.100 50.600 75.200 ;
        RECT 54.200 75.100 54.600 75.200 ;
        RECT 50.200 74.800 54.600 75.100 ;
        RECT 62.200 75.100 62.600 75.200 ;
        RECT 66.200 75.100 66.600 75.200 ;
        RECT 71.800 75.100 72.200 75.200 ;
        RECT 62.200 74.800 72.200 75.100 ;
        RECT 75.000 75.100 75.400 75.200 ;
        RECT 80.600 75.100 81.000 75.200 ;
        RECT 75.000 74.800 81.000 75.100 ;
        RECT 99.000 74.800 99.400 75.200 ;
        RECT 104.600 75.100 105.000 75.200 ;
        RECT 105.400 75.100 105.800 75.200 ;
        RECT 104.600 74.800 105.800 75.100 ;
        RECT 139.000 74.800 139.400 75.200 ;
        RECT 142.200 75.100 142.600 75.200 ;
        RECT 145.400 75.100 145.700 75.800 ;
        RECT 142.200 74.800 145.700 75.100 ;
        RECT 7.800 74.100 8.200 74.200 ;
        RECT 13.400 74.100 13.800 74.200 ;
        RECT 15.000 74.100 15.400 74.200 ;
        RECT 7.800 73.800 15.400 74.100 ;
        RECT 18.200 73.800 18.600 74.200 ;
        RECT 19.000 74.100 19.400 74.200 ;
        RECT 23.800 74.100 24.200 74.200 ;
        RECT 29.400 74.100 29.800 74.200 ;
        RECT 19.000 73.800 22.500 74.100 ;
        RECT 23.800 73.800 29.800 74.100 ;
        RECT 33.400 74.100 33.800 74.200 ;
        RECT 39.000 74.100 39.400 74.200 ;
        RECT 33.400 73.800 39.400 74.100 ;
        RECT 52.600 73.800 53.000 74.200 ;
        RECT 60.600 74.100 61.000 74.200 ;
        RECT 61.400 74.100 61.800 74.200 ;
        RECT 60.600 73.800 61.800 74.100 ;
        RECT 72.600 74.100 73.000 74.200 ;
        RECT 90.200 74.100 90.600 74.200 ;
        RECT 108.600 74.100 109.000 74.200 ;
        RECT 72.600 73.800 109.000 74.100 ;
        RECT 112.600 74.100 113.000 74.200 ;
        RECT 113.400 74.100 113.800 74.200 ;
        RECT 119.000 74.100 119.400 74.200 ;
        RECT 112.600 73.800 119.400 74.100 ;
        RECT 121.400 74.100 121.800 74.200 ;
        RECT 123.000 74.100 123.400 74.200 ;
        RECT 125.400 74.100 125.800 74.200 ;
        RECT 121.400 73.800 125.800 74.100 ;
        RECT 130.200 74.100 130.600 74.200 ;
        RECT 132.600 74.100 133.000 74.200 ;
        RECT 130.200 73.800 133.000 74.100 ;
        RECT 135.800 74.100 136.200 74.200 ;
        RECT 143.000 74.100 143.400 74.200 ;
        RECT 135.800 73.800 143.400 74.100 ;
        RECT 11.800 73.200 12.100 73.800 ;
        RECT 18.200 73.200 18.500 73.800 ;
        RECT 22.200 73.200 22.500 73.800 ;
        RECT 52.600 73.200 52.900 73.800 ;
        RECT 8.600 73.100 9.000 73.200 ;
        RECT 9.400 73.100 9.800 73.200 ;
        RECT 8.600 72.800 9.800 73.100 ;
        RECT 11.800 72.800 12.200 73.200 ;
        RECT 16.600 73.100 17.000 73.200 ;
        RECT 17.400 73.100 17.800 73.200 ;
        RECT 16.600 72.800 17.800 73.100 ;
        RECT 18.200 72.800 18.600 73.200 ;
        RECT 22.200 72.800 22.600 73.200 ;
        RECT 25.400 73.100 25.800 73.200 ;
        RECT 27.000 73.100 27.400 73.200 ;
        RECT 25.400 72.800 27.400 73.100 ;
        RECT 34.200 73.100 34.600 73.200 ;
        RECT 42.200 73.100 42.600 73.200 ;
        RECT 43.800 73.100 44.200 73.200 ;
        RECT 34.200 72.800 44.200 73.100 ;
        RECT 45.400 72.800 45.800 73.200 ;
        RECT 52.600 72.800 53.000 73.200 ;
        RECT 59.000 73.100 59.400 73.200 ;
        RECT 81.400 73.100 81.800 73.200 ;
        RECT 59.000 72.800 81.800 73.100 ;
        RECT 83.800 73.100 84.200 73.200 ;
        RECT 84.600 73.100 85.000 73.200 ;
        RECT 83.800 72.800 85.000 73.100 ;
        RECT 91.800 72.800 92.200 73.200 ;
        RECT 94.200 73.100 94.600 73.200 ;
        RECT 100.600 73.100 101.000 73.200 ;
        RECT 94.200 72.800 101.000 73.100 ;
        RECT 101.400 73.100 101.800 73.200 ;
        RECT 104.600 73.100 105.000 73.200 ;
        RECT 101.400 72.800 105.000 73.100 ;
        RECT 111.800 73.100 112.200 73.200 ;
        RECT 115.000 73.100 115.400 73.200 ;
        RECT 111.800 72.800 115.400 73.100 ;
        RECT 120.600 73.100 121.000 73.200 ;
        RECT 122.200 73.100 122.600 73.200 ;
        RECT 120.600 72.800 122.600 73.100 ;
        RECT 141.400 72.800 141.800 73.200 ;
        RECT 45.400 72.200 45.700 72.800 ;
        RECT 21.400 72.100 21.800 72.200 ;
        RECT 25.400 72.100 25.800 72.200 ;
        RECT 35.000 72.100 35.400 72.200 ;
        RECT 21.400 71.800 35.400 72.100 ;
        RECT 36.600 72.100 37.000 72.200 ;
        RECT 44.600 72.100 45.000 72.200 ;
        RECT 36.600 71.800 45.000 72.100 ;
        RECT 45.400 71.800 45.800 72.200 ;
        RECT 60.600 72.100 61.000 72.200 ;
        RECT 68.600 72.100 69.000 72.200 ;
        RECT 60.600 71.800 69.000 72.100 ;
        RECT 69.400 72.100 69.800 72.200 ;
        RECT 70.200 72.100 70.600 72.200 ;
        RECT 69.400 71.800 70.600 72.100 ;
        RECT 71.800 72.100 72.200 72.200 ;
        RECT 79.800 72.100 80.200 72.200 ;
        RECT 83.000 72.100 83.400 72.200 ;
        RECT 86.200 72.100 86.600 72.200 ;
        RECT 71.800 71.800 86.600 72.100 ;
        RECT 91.800 72.100 92.100 72.800 ;
        RECT 141.400 72.200 141.700 72.800 ;
        RECT 95.000 72.100 95.400 72.200 ;
        RECT 91.800 71.800 95.400 72.100 ;
        RECT 95.800 72.100 96.200 72.200 ;
        RECT 104.600 72.100 105.000 72.200 ;
        RECT 95.800 71.800 105.000 72.100 ;
        RECT 105.400 72.100 105.800 72.200 ;
        RECT 119.800 72.100 120.200 72.200 ;
        RECT 126.200 72.100 126.600 72.200 ;
        RECT 105.400 71.800 126.600 72.100 ;
        RECT 141.400 71.800 141.800 72.200 ;
        RECT 15.000 71.100 15.400 71.200 ;
        RECT 26.200 71.100 26.600 71.200 ;
        RECT 15.000 70.800 26.600 71.100 ;
        RECT 39.000 71.100 39.400 71.200 ;
        RECT 39.800 71.100 40.200 71.200 ;
        RECT 39.000 70.800 40.200 71.100 ;
        RECT 55.000 71.100 55.400 71.200 ;
        RECT 57.400 71.100 57.800 71.200 ;
        RECT 55.000 70.800 57.800 71.100 ;
        RECT 65.400 71.100 65.800 71.200 ;
        RECT 77.400 71.100 77.800 71.200 ;
        RECT 65.400 70.800 77.800 71.100 ;
        RECT 87.000 71.100 87.400 71.200 ;
        RECT 98.200 71.100 98.600 71.200 ;
        RECT 87.000 70.800 98.600 71.100 ;
        RECT 103.000 71.100 103.400 71.200 ;
        RECT 105.400 71.100 105.800 71.200 ;
        RECT 103.000 70.800 105.800 71.100 ;
        RECT 107.000 71.100 107.400 71.200 ;
        RECT 111.000 71.100 111.400 71.200 ;
        RECT 130.200 71.100 130.600 71.200 ;
        RECT 147.000 71.100 147.400 71.200 ;
        RECT 107.000 70.800 147.400 71.100 ;
        RECT 27.800 70.100 28.200 70.200 ;
        RECT 34.200 70.100 34.600 70.200 ;
        RECT 27.800 69.800 34.600 70.100 ;
        RECT 35.000 70.100 35.400 70.200 ;
        RECT 36.600 70.100 37.000 70.200 ;
        RECT 35.000 69.800 37.000 70.100 ;
        RECT 38.200 70.100 38.600 70.200 ;
        RECT 114.200 70.100 114.600 70.200 ;
        RECT 115.000 70.100 115.400 70.200 ;
        RECT 38.200 69.800 99.300 70.100 ;
        RECT 114.200 69.800 115.400 70.100 ;
        RECT 116.600 70.100 117.000 70.200 ;
        RECT 125.400 70.100 125.800 70.200 ;
        RECT 116.600 69.800 125.800 70.100 ;
        RECT 140.600 70.100 141.000 70.200 ;
        RECT 143.800 70.100 144.200 70.200 ;
        RECT 140.600 69.800 144.200 70.100 ;
        RECT 0.600 69.100 1.000 69.200 ;
        RECT 20.600 69.100 21.000 69.200 ;
        RECT 22.200 69.100 22.600 69.200 ;
        RECT 30.200 69.100 30.600 69.200 ;
        RECT 31.000 69.100 31.400 69.200 ;
        RECT 35.800 69.100 36.200 69.200 ;
        RECT 0.600 68.800 4.900 69.100 ;
        RECT 20.600 68.800 36.200 69.100 ;
        RECT 39.800 69.100 40.200 69.200 ;
        RECT 55.800 69.100 56.200 69.200 ;
        RECT 61.400 69.100 61.800 69.200 ;
        RECT 39.800 68.800 45.700 69.100 ;
        RECT 55.800 68.800 61.800 69.100 ;
        RECT 66.200 69.100 66.600 69.200 ;
        RECT 67.800 69.100 68.200 69.200 ;
        RECT 66.200 68.800 68.200 69.100 ;
        RECT 68.600 69.100 69.000 69.200 ;
        RECT 75.000 69.100 75.400 69.200 ;
        RECT 81.400 69.100 81.800 69.200 ;
        RECT 68.600 68.800 81.800 69.100 ;
        RECT 99.000 69.100 99.300 69.800 ;
        RECT 128.600 69.100 129.000 69.200 ;
        RECT 99.000 68.800 129.000 69.100 ;
        RECT 133.400 69.100 133.800 69.200 ;
        RECT 146.200 69.100 146.600 69.200 ;
        RECT 133.400 68.800 146.600 69.100 ;
        RECT 4.600 68.200 4.900 68.800 ;
        RECT 45.400 68.200 45.700 68.800 ;
        RECT 4.600 67.800 5.000 68.200 ;
        RECT 21.400 68.100 21.800 68.200 ;
        RECT 24.600 68.100 25.000 68.200 ;
        RECT 28.600 68.100 29.000 68.200 ;
        RECT 38.200 68.100 38.600 68.200 ;
        RECT 21.400 67.800 38.600 68.100 ;
        RECT 45.400 67.800 45.800 68.200 ;
        RECT 58.200 68.100 58.600 68.200 ;
        RECT 63.000 68.100 63.400 68.200 ;
        RECT 58.200 67.800 63.400 68.100 ;
        RECT 64.600 68.100 65.000 68.200 ;
        RECT 69.400 68.100 69.800 68.200 ;
        RECT 64.600 67.800 69.800 68.100 ;
        RECT 70.200 68.100 70.600 68.200 ;
        RECT 71.000 68.100 71.400 68.200 ;
        RECT 111.800 68.100 112.200 68.200 ;
        RECT 70.200 67.800 71.400 68.100 ;
        RECT 98.200 67.800 112.200 68.100 ;
        RECT 115.800 68.100 116.200 68.200 ;
        RECT 117.400 68.100 117.800 68.200 ;
        RECT 115.800 67.800 117.800 68.100 ;
        RECT 118.200 68.100 118.600 68.200 ;
        RECT 123.000 68.100 123.400 68.200 ;
        RECT 118.200 67.800 123.400 68.100 ;
        RECT 123.800 68.100 124.200 68.200 ;
        RECT 126.200 68.100 126.600 68.200 ;
        RECT 139.000 68.100 139.400 68.200 ;
        RECT 123.800 67.800 126.600 68.100 ;
        RECT 131.800 67.800 139.400 68.100 ;
        RECT 98.200 67.200 98.500 67.800 ;
        RECT 131.800 67.200 132.100 67.800 ;
        RECT 8.600 67.100 9.000 67.200 ;
        RECT 11.000 67.100 11.400 67.200 ;
        RECT 94.200 67.100 94.600 67.200 ;
        RECT 8.600 66.800 11.400 67.100 ;
        RECT 84.600 66.800 94.600 67.100 ;
        RECT 96.600 66.800 97.000 67.200 ;
        RECT 98.200 66.800 98.600 67.200 ;
        RECT 103.800 67.100 104.200 67.200 ;
        RECT 104.600 67.100 105.000 67.200 ;
        RECT 103.800 66.800 105.000 67.100 ;
        RECT 112.600 67.100 113.000 67.200 ;
        RECT 120.600 67.100 121.000 67.200 ;
        RECT 112.600 66.800 121.000 67.100 ;
        RECT 123.000 66.800 123.400 67.200 ;
        RECT 125.400 67.100 125.800 67.200 ;
        RECT 127.000 67.100 127.400 67.200 ;
        RECT 125.400 66.800 127.400 67.100 ;
        RECT 131.800 66.800 132.200 67.200 ;
        RECT 132.600 67.100 133.000 67.200 ;
        RECT 136.600 67.100 137.000 67.200 ;
        RECT 132.600 66.800 137.000 67.100 ;
        RECT 5.400 66.100 5.800 66.200 ;
        RECT 9.400 66.100 9.800 66.200 ;
        RECT 5.400 65.800 9.800 66.100 ;
        RECT 14.200 66.100 14.600 66.200 ;
        RECT 15.800 66.100 16.200 66.200 ;
        RECT 14.200 65.800 16.200 66.100 ;
        RECT 19.800 66.100 20.200 66.200 ;
        RECT 23.800 66.100 24.200 66.200 ;
        RECT 19.800 65.800 24.200 66.100 ;
        RECT 27.000 65.800 27.400 66.200 ;
        RECT 63.800 66.100 64.200 66.200 ;
        RECT 74.200 66.100 74.600 66.200 ;
        RECT 63.800 65.800 74.600 66.100 ;
        RECT 78.200 66.100 78.600 66.200 ;
        RECT 84.600 66.100 84.900 66.800 ;
        RECT 78.200 65.800 84.900 66.100 ;
        RECT 91.000 66.100 91.400 66.200 ;
        RECT 96.600 66.100 96.900 66.800 ;
        RECT 123.000 66.200 123.300 66.800 ;
        RECT 91.000 65.800 96.900 66.100 ;
        RECT 106.200 66.100 106.600 66.200 ;
        RECT 108.600 66.100 109.000 66.200 ;
        RECT 106.200 65.800 109.000 66.100 ;
        RECT 111.800 66.100 112.200 66.200 ;
        RECT 115.800 66.100 116.200 66.200 ;
        RECT 119.000 66.100 119.400 66.200 ;
        RECT 111.800 65.800 119.400 66.100 ;
        RECT 123.000 65.800 123.400 66.200 ;
        RECT 127.800 66.100 128.200 66.200 ;
        RECT 130.200 66.100 130.600 66.200 ;
        RECT 135.000 66.100 135.400 66.200 ;
        RECT 127.800 65.800 135.400 66.100 ;
        RECT 27.000 65.200 27.300 65.800 ;
        RECT 0.600 65.100 1.000 65.200 ;
        RECT 2.200 65.100 2.600 65.200 ;
        RECT 6.200 65.100 6.600 65.200 ;
        RECT 0.600 64.800 6.600 65.100 ;
        RECT 8.600 65.100 9.000 65.200 ;
        RECT 10.200 65.100 10.600 65.200 ;
        RECT 8.600 64.800 10.600 65.100 ;
        RECT 11.800 65.100 12.200 65.200 ;
        RECT 17.400 65.100 17.800 65.200 ;
        RECT 11.800 64.800 17.800 65.100 ;
        RECT 27.000 64.800 27.400 65.200 ;
        RECT 39.800 65.100 40.200 65.200 ;
        RECT 52.600 65.100 53.000 65.200 ;
        RECT 39.800 64.800 53.000 65.100 ;
        RECT 88.600 65.100 89.000 65.200 ;
        RECT 99.000 65.100 99.400 65.200 ;
        RECT 88.600 64.800 99.400 65.100 ;
        RECT 104.600 65.100 105.000 65.200 ;
        RECT 112.600 65.100 113.000 65.200 ;
        RECT 104.600 64.800 113.000 65.100 ;
        RECT 116.600 65.100 117.000 65.200 ;
        RECT 118.200 65.100 118.600 65.200 ;
        RECT 116.600 64.800 118.600 65.100 ;
        RECT 124.600 65.100 125.000 65.200 ;
        RECT 127.800 65.100 128.200 65.200 ;
        RECT 128.600 65.100 129.000 65.200 ;
        RECT 124.600 64.800 129.000 65.100 ;
        RECT 137.400 64.800 140.900 65.100 ;
        RECT 15.800 64.200 16.100 64.800 ;
        RECT 137.400 64.200 137.700 64.800 ;
        RECT 140.600 64.200 140.900 64.800 ;
        RECT 8.600 64.100 9.000 64.200 ;
        RECT 14.200 64.100 14.600 64.200 ;
        RECT 8.600 63.800 14.600 64.100 ;
        RECT 15.800 63.800 16.200 64.200 ;
        RECT 16.600 64.100 17.000 64.200 ;
        RECT 19.000 64.100 19.400 64.200 ;
        RECT 16.600 63.800 19.400 64.100 ;
        RECT 60.600 64.100 61.000 64.200 ;
        RECT 68.600 64.100 69.000 64.200 ;
        RECT 60.600 63.800 69.000 64.100 ;
        RECT 90.200 64.100 90.600 64.200 ;
        RECT 101.400 64.100 101.800 64.200 ;
        RECT 90.200 63.800 101.800 64.100 ;
        RECT 107.800 64.100 108.200 64.200 ;
        RECT 125.400 64.100 125.800 64.200 ;
        RECT 107.800 63.800 125.800 64.100 ;
        RECT 132.600 64.100 133.000 64.200 ;
        RECT 133.400 64.100 133.800 64.200 ;
        RECT 132.600 63.800 133.800 64.100 ;
        RECT 137.400 63.800 137.800 64.200 ;
        RECT 140.600 63.800 141.000 64.200 ;
        RECT 143.800 64.100 144.200 64.200 ;
        RECT 147.000 64.100 147.400 64.200 ;
        RECT 143.800 63.800 147.400 64.100 ;
        RECT 7.800 63.100 8.200 63.200 ;
        RECT 26.200 63.100 26.600 63.200 ;
        RECT 7.800 62.800 26.600 63.100 ;
        RECT 42.200 63.100 42.600 63.200 ;
        RECT 55.800 63.100 56.200 63.200 ;
        RECT 42.200 62.800 56.200 63.100 ;
        RECT 63.800 63.100 64.200 63.200 ;
        RECT 72.600 63.100 73.000 63.200 ;
        RECT 63.800 62.800 73.000 63.100 ;
        RECT 76.600 63.100 77.000 63.200 ;
        RECT 92.600 63.100 93.000 63.200 ;
        RECT 76.600 62.800 93.000 63.100 ;
        RECT 99.800 63.100 100.200 63.200 ;
        RECT 142.200 63.100 142.600 63.200 ;
        RECT 99.800 62.800 142.600 63.100 ;
        RECT 44.600 62.100 45.000 62.200 ;
        RECT 76.600 62.100 77.000 62.200 ;
        RECT 44.600 61.800 77.000 62.100 ;
        RECT 79.800 62.100 80.200 62.200 ;
        RECT 82.200 62.100 82.600 62.200 ;
        RECT 93.400 62.100 93.800 62.200 ;
        RECT 111.800 62.100 112.200 62.200 ;
        RECT 120.600 62.100 121.000 62.200 ;
        RECT 79.800 61.800 82.600 62.100 ;
        RECT 92.600 61.800 121.000 62.100 ;
        RECT 123.000 62.100 123.400 62.200 ;
        RECT 132.600 62.100 133.000 62.200 ;
        RECT 123.000 61.800 133.000 62.100 ;
        RECT 135.800 62.100 136.200 62.200 ;
        RECT 145.400 62.100 145.800 62.200 ;
        RECT 135.800 61.800 145.800 62.100 ;
        RECT 14.200 61.100 14.600 61.200 ;
        RECT 21.400 61.100 21.800 61.200 ;
        RECT 14.200 60.800 21.800 61.100 ;
        RECT 55.000 61.100 55.400 61.200 ;
        RECT 60.600 61.100 61.000 61.200 ;
        RECT 75.000 61.100 75.400 61.200 ;
        RECT 111.800 61.100 112.200 61.200 ;
        RECT 55.000 60.800 74.500 61.100 ;
        RECT 75.000 60.800 112.200 61.100 ;
        RECT 15.800 60.100 16.200 60.200 ;
        RECT 35.000 60.100 35.400 60.200 ;
        RECT 15.800 59.800 35.400 60.100 ;
        RECT 74.200 60.100 74.500 60.800 ;
        RECT 81.400 60.100 81.800 60.200 ;
        RECT 84.600 60.100 85.000 60.200 ;
        RECT 91.000 60.100 91.400 60.200 ;
        RECT 74.200 59.800 91.400 60.100 ;
        RECT 101.400 60.100 101.800 60.200 ;
        RECT 124.600 60.100 125.000 60.200 ;
        RECT 101.400 59.800 125.000 60.100 ;
        RECT 24.600 58.800 25.000 59.200 ;
        RECT 45.400 59.100 45.800 59.200 ;
        RECT 48.600 59.100 49.000 59.200 ;
        RECT 45.400 58.800 49.000 59.100 ;
        RECT 50.200 59.100 50.600 59.200 ;
        RECT 58.200 59.100 58.600 59.200 ;
        RECT 50.200 58.800 58.600 59.100 ;
        RECT 98.200 59.100 98.600 59.200 ;
        RECT 143.800 59.100 144.200 59.200 ;
        RECT 98.200 58.800 144.200 59.100 ;
        RECT 5.400 57.800 5.800 58.200 ;
        RECT 19.800 58.100 20.200 58.200 ;
        RECT 24.600 58.100 24.900 58.800 ;
        RECT 19.800 57.800 24.900 58.100 ;
        RECT 54.200 58.100 54.600 58.200 ;
        RECT 63.000 58.100 63.400 58.200 ;
        RECT 71.800 58.100 72.200 58.200 ;
        RECT 54.200 57.800 72.200 58.100 ;
        RECT 79.000 57.800 79.400 58.200 ;
        RECT 80.600 58.100 81.000 58.200 ;
        RECT 89.400 58.100 89.800 58.200 ;
        RECT 100.600 58.100 101.000 58.200 ;
        RECT 80.600 57.800 101.000 58.100 ;
        RECT 105.400 58.100 105.800 58.200 ;
        RECT 124.600 58.100 125.000 58.200 ;
        RECT 132.600 58.100 133.000 58.200 ;
        RECT 105.400 57.800 133.000 58.100 ;
        RECT 135.000 57.800 135.400 58.200 ;
        RECT 4.600 57.100 5.000 57.200 ;
        RECT 5.400 57.100 5.700 57.800 ;
        RECT 4.600 56.800 5.700 57.100 ;
        RECT 10.200 57.100 10.600 57.200 ;
        RECT 11.000 57.100 11.400 57.200 ;
        RECT 10.200 56.800 11.400 57.100 ;
        RECT 23.000 57.100 23.400 57.200 ;
        RECT 25.400 57.100 25.800 57.200 ;
        RECT 23.000 56.800 25.800 57.100 ;
        RECT 32.600 57.100 33.000 57.200 ;
        RECT 36.600 57.100 37.000 57.200 ;
        RECT 32.600 56.800 37.000 57.100 ;
        RECT 37.400 57.100 37.800 57.200 ;
        RECT 69.400 57.100 69.800 57.200 ;
        RECT 37.400 56.800 69.800 57.100 ;
        RECT 79.000 57.100 79.300 57.800 ;
        RECT 92.600 57.100 93.000 57.200 ;
        RECT 79.000 56.800 93.000 57.100 ;
        RECT 101.400 56.800 101.800 57.200 ;
        RECT 104.600 57.100 105.000 57.200 ;
        RECT 111.000 57.100 111.400 57.200 ;
        RECT 104.600 56.800 111.400 57.100 ;
        RECT 113.400 56.800 113.800 57.200 ;
        RECT 115.000 57.100 115.400 57.200 ;
        RECT 126.200 57.100 126.600 57.200 ;
        RECT 135.000 57.100 135.300 57.800 ;
        RECT 115.000 56.800 126.600 57.100 ;
        RECT 130.200 56.800 135.300 57.100 ;
        RECT 15.000 56.100 15.400 56.200 ;
        RECT 17.400 56.100 17.800 56.200 ;
        RECT 15.000 55.800 17.800 56.100 ;
        RECT 19.000 56.100 19.400 56.200 ;
        RECT 31.800 56.100 32.200 56.200 ;
        RECT 19.000 55.800 32.200 56.100 ;
        RECT 67.000 56.100 67.400 56.200 ;
        RECT 75.000 56.100 75.400 56.200 ;
        RECT 67.000 55.800 75.400 56.100 ;
        RECT 75.800 56.100 76.200 56.200 ;
        RECT 76.600 56.100 77.000 56.200 ;
        RECT 75.800 55.800 77.000 56.100 ;
        RECT 81.400 56.100 81.800 56.200 ;
        RECT 87.000 56.100 87.400 56.200 ;
        RECT 81.400 55.800 87.400 56.100 ;
        RECT 98.200 56.100 98.600 56.200 ;
        RECT 101.400 56.100 101.700 56.800 ;
        RECT 113.400 56.200 113.700 56.800 ;
        RECT 130.200 56.200 130.500 56.800 ;
        RECT 98.200 55.800 101.700 56.100 ;
        RECT 106.200 56.100 106.600 56.200 ;
        RECT 108.600 56.100 109.000 56.200 ;
        RECT 106.200 55.800 109.000 56.100 ;
        RECT 110.200 56.100 110.600 56.200 ;
        RECT 111.000 56.100 111.400 56.200 ;
        RECT 110.200 55.800 111.400 56.100 ;
        RECT 113.400 55.800 113.800 56.200 ;
        RECT 119.000 56.100 119.400 56.200 ;
        RECT 119.000 55.800 122.500 56.100 ;
        RECT 130.200 55.800 130.600 56.200 ;
        RECT 133.400 55.800 133.800 56.200 ;
        RECT 122.200 55.200 122.500 55.800 ;
        RECT 133.400 55.200 133.700 55.800 ;
        RECT 3.800 55.100 4.200 55.200 ;
        RECT 10.200 55.100 10.600 55.200 ;
        RECT 3.800 54.800 10.600 55.100 ;
        RECT 11.000 55.100 11.400 55.200 ;
        RECT 12.600 55.100 13.000 55.200 ;
        RECT 11.000 54.800 13.000 55.100 ;
        RECT 22.200 55.100 22.600 55.200 ;
        RECT 26.200 55.100 26.600 55.200 ;
        RECT 22.200 54.800 26.600 55.100 ;
        RECT 29.400 55.100 29.800 55.200 ;
        RECT 31.800 55.100 32.200 55.200 ;
        RECT 35.800 55.100 36.200 55.200 ;
        RECT 29.400 54.800 36.200 55.100 ;
        RECT 39.000 54.800 39.400 55.200 ;
        RECT 40.600 55.100 41.000 55.200 ;
        RECT 41.400 55.100 41.800 55.200 ;
        RECT 40.600 54.800 41.800 55.100 ;
        RECT 42.200 55.100 42.600 55.200 ;
        RECT 45.400 55.100 45.800 55.200 ;
        RECT 42.200 54.800 45.800 55.100 ;
        RECT 53.400 55.100 53.800 55.200 ;
        RECT 54.200 55.100 54.600 55.200 ;
        RECT 53.400 54.800 54.600 55.100 ;
        RECT 60.600 55.100 61.000 55.200 ;
        RECT 64.600 55.100 65.000 55.200 ;
        RECT 67.000 55.100 67.400 55.200 ;
        RECT 60.600 54.800 67.400 55.100 ;
        RECT 71.800 55.100 72.200 55.200 ;
        RECT 72.600 55.100 73.000 55.200 ;
        RECT 79.800 55.100 80.200 55.200 ;
        RECT 71.800 54.800 80.200 55.100 ;
        RECT 91.000 55.100 91.400 55.200 ;
        RECT 93.400 55.100 93.800 55.200 ;
        RECT 91.000 54.800 93.800 55.100 ;
        RECT 97.400 55.100 97.800 55.200 ;
        RECT 99.800 55.100 100.200 55.200 ;
        RECT 97.400 54.800 100.200 55.100 ;
        RECT 101.400 55.100 101.800 55.200 ;
        RECT 106.200 55.100 106.600 55.200 ;
        RECT 107.800 55.100 108.200 55.200 ;
        RECT 101.400 54.800 108.200 55.100 ;
        RECT 115.000 55.100 115.400 55.200 ;
        RECT 115.800 55.100 116.200 55.200 ;
        RECT 115.000 54.800 116.200 55.100 ;
        RECT 120.600 55.100 121.000 55.200 ;
        RECT 121.400 55.100 121.800 55.200 ;
        RECT 120.600 54.800 121.800 55.100 ;
        RECT 122.200 54.800 122.600 55.200 ;
        RECT 123.000 55.100 123.400 55.200 ;
        RECT 123.800 55.100 124.200 55.200 ;
        RECT 123.000 54.800 124.200 55.100 ;
        RECT 133.400 54.800 133.800 55.200 ;
        RECT 145.400 55.100 145.800 55.200 ;
        RECT 147.000 55.100 147.400 55.200 ;
        RECT 145.400 54.800 147.400 55.100 ;
        RECT 148.600 55.100 149.000 55.200 ;
        RECT 149.400 55.100 149.800 55.200 ;
        RECT 148.600 54.800 149.800 55.100 ;
        RECT 15.000 54.100 15.400 54.200 ;
        RECT 17.400 54.100 17.800 54.200 ;
        RECT 15.000 53.800 17.800 54.100 ;
        RECT 23.800 54.100 24.200 54.200 ;
        RECT 24.600 54.100 25.000 54.200 ;
        RECT 31.000 54.100 31.400 54.200 ;
        RECT 39.000 54.100 39.300 54.800 ;
        RECT 23.800 53.800 39.300 54.100 ;
        RECT 60.600 53.800 61.000 54.200 ;
        RECT 67.000 54.100 67.400 54.200 ;
        RECT 68.600 54.100 69.000 54.200 ;
        RECT 67.000 53.800 69.000 54.100 ;
        RECT 71.000 54.100 71.400 54.200 ;
        RECT 79.800 54.100 80.200 54.200 ;
        RECT 71.000 53.800 80.200 54.100 ;
        RECT 88.600 54.100 89.000 54.200 ;
        RECT 89.400 54.100 89.800 54.200 ;
        RECT 88.600 53.800 89.800 54.100 ;
        RECT 95.000 54.100 95.400 54.200 ;
        RECT 101.400 54.100 101.800 54.200 ;
        RECT 95.000 53.800 101.800 54.100 ;
        RECT 103.800 53.800 104.200 54.200 ;
        RECT 104.600 54.100 105.000 54.200 ;
        RECT 108.600 54.100 109.000 54.200 ;
        RECT 104.600 53.800 109.000 54.100 ;
        RECT 124.600 54.100 125.000 54.200 ;
        RECT 126.200 54.100 126.600 54.200 ;
        RECT 124.600 53.800 126.600 54.100 ;
        RECT 137.400 54.100 137.800 54.200 ;
        RECT 143.000 54.100 143.400 54.200 ;
        RECT 137.400 53.800 143.400 54.100 ;
        RECT 148.600 53.800 149.000 54.200 ;
        RECT 60.600 53.200 60.900 53.800 ;
        RECT 28.600 53.100 29.000 53.200 ;
        RECT 34.200 53.100 34.600 53.200 ;
        RECT 51.000 53.100 51.400 53.200 ;
        RECT 52.600 53.100 53.000 53.200 ;
        RECT 53.400 53.100 53.800 53.200 ;
        RECT 28.600 52.800 46.500 53.100 ;
        RECT 51.000 52.800 53.800 53.100 ;
        RECT 60.600 52.800 61.000 53.200 ;
        RECT 87.800 53.100 88.200 53.200 ;
        RECT 91.800 53.100 92.200 53.200 ;
        RECT 93.400 53.100 93.800 53.200 ;
        RECT 87.800 52.800 93.800 53.100 ;
        RECT 102.200 53.100 102.600 53.200 ;
        RECT 103.000 53.100 103.400 53.200 ;
        RECT 102.200 52.800 103.400 53.100 ;
        RECT 103.800 53.100 104.100 53.800 ;
        RECT 104.600 53.100 105.000 53.200 ;
        RECT 103.800 52.800 105.000 53.100 ;
        RECT 107.800 53.100 108.200 53.200 ;
        RECT 109.400 53.100 109.800 53.200 ;
        RECT 119.000 53.100 119.400 53.200 ;
        RECT 143.000 53.100 143.400 53.200 ;
        RECT 107.800 52.800 119.400 53.100 ;
        RECT 125.400 52.800 143.400 53.100 ;
        RECT 147.000 53.100 147.400 53.200 ;
        RECT 148.600 53.100 148.900 53.800 ;
        RECT 147.000 52.800 148.900 53.100 ;
        RECT 46.200 52.200 46.500 52.800 ;
        RECT 125.400 52.200 125.700 52.800 ;
        RECT 0.600 52.100 1.000 52.200 ;
        RECT 15.800 52.100 16.200 52.200 ;
        RECT 0.600 51.800 16.200 52.100 ;
        RECT 17.400 52.100 17.800 52.200 ;
        RECT 27.800 52.100 28.200 52.200 ;
        RECT 17.400 51.800 28.200 52.100 ;
        RECT 29.400 52.100 29.800 52.200 ;
        RECT 32.600 52.100 33.000 52.200 ;
        RECT 37.400 52.100 37.800 52.200 ;
        RECT 29.400 51.800 37.800 52.100 ;
        RECT 46.200 51.800 46.600 52.200 ;
        RECT 51.800 52.100 52.200 52.200 ;
        RECT 55.000 52.100 55.400 52.200 ;
        RECT 51.800 51.800 55.400 52.100 ;
        RECT 76.600 52.100 77.000 52.200 ;
        RECT 77.400 52.100 77.800 52.200 ;
        RECT 76.600 51.800 77.800 52.100 ;
        RECT 82.200 52.100 82.600 52.200 ;
        RECT 85.400 52.100 85.800 52.200 ;
        RECT 82.200 51.800 85.800 52.100 ;
        RECT 107.000 52.100 107.400 52.200 ;
        RECT 107.800 52.100 108.200 52.200 ;
        RECT 107.000 51.800 108.200 52.100 ;
        RECT 125.400 51.800 125.800 52.200 ;
        RECT 126.200 52.100 126.600 52.200 ;
        RECT 129.400 52.100 129.800 52.200 ;
        RECT 136.600 52.100 137.000 52.200 ;
        RECT 126.200 51.800 137.000 52.100 ;
        RECT 142.200 52.100 142.600 52.200 ;
        RECT 147.000 52.100 147.300 52.800 ;
        RECT 142.200 51.800 147.300 52.100 ;
        RECT 13.400 51.100 13.800 51.200 ;
        RECT 25.400 51.100 25.800 51.200 ;
        RECT 13.400 50.800 25.800 51.100 ;
        RECT 69.400 51.100 69.800 51.200 ;
        RECT 70.200 51.100 70.600 51.200 ;
        RECT 69.400 50.800 70.600 51.100 ;
        RECT 71.800 51.100 72.200 51.200 ;
        RECT 79.000 51.100 79.400 51.200 ;
        RECT 71.800 50.800 79.400 51.100 ;
        RECT 83.800 51.100 84.200 51.200 ;
        RECT 98.200 51.100 98.600 51.200 ;
        RECT 83.800 50.800 98.600 51.100 ;
        RECT 105.400 51.100 105.800 51.200 ;
        RECT 113.400 51.100 113.800 51.200 ;
        RECT 105.400 50.800 113.800 51.100 ;
        RECT 119.000 51.100 119.400 51.200 ;
        RECT 141.400 51.100 141.800 51.200 ;
        RECT 119.000 50.800 141.800 51.100 ;
        RECT 149.400 51.100 149.800 51.200 ;
        RECT 150.200 51.100 150.600 51.200 ;
        RECT 149.400 50.800 150.600 51.100 ;
        RECT 16.600 50.100 17.000 50.200 ;
        RECT 23.800 50.100 24.200 50.200 ;
        RECT 16.600 49.800 24.200 50.100 ;
        RECT 47.000 50.100 47.400 50.200 ;
        RECT 54.200 50.100 54.600 50.200 ;
        RECT 47.000 49.800 54.600 50.100 ;
        RECT 55.000 50.100 55.400 50.200 ;
        RECT 61.400 50.100 61.800 50.200 ;
        RECT 55.000 49.800 61.800 50.100 ;
        RECT 63.000 50.100 63.400 50.200 ;
        RECT 83.800 50.100 84.200 50.200 ;
        RECT 63.000 49.800 84.200 50.100 ;
        RECT 95.800 50.100 96.200 50.200 ;
        RECT 97.400 50.100 97.800 50.200 ;
        RECT 95.800 49.800 97.800 50.100 ;
        RECT 124.600 50.100 125.000 50.200 ;
        RECT 138.200 50.100 138.600 50.200 ;
        RECT 124.600 49.800 138.600 50.100 ;
        RECT 147.800 50.100 148.200 50.200 ;
        RECT 149.400 50.100 149.800 50.200 ;
        RECT 147.800 49.800 149.800 50.100 ;
        RECT 7.000 49.100 7.400 49.200 ;
        RECT 9.400 49.100 9.800 49.200 ;
        RECT 18.200 49.100 18.600 49.200 ;
        RECT 67.800 49.100 68.200 49.200 ;
        RECT 7.000 48.800 68.200 49.100 ;
        RECT 69.400 49.100 69.800 49.200 ;
        RECT 77.400 49.100 77.800 49.200 ;
        RECT 69.400 48.800 77.800 49.100 ;
        RECT 82.200 49.100 82.600 49.200 ;
        RECT 97.400 49.100 97.800 49.200 ;
        RECT 82.200 48.800 97.800 49.100 ;
        RECT 99.000 49.100 99.400 49.200 ;
        RECT 105.400 49.100 105.800 49.200 ;
        RECT 99.000 48.800 105.800 49.100 ;
        RECT 111.800 48.800 112.200 49.200 ;
        RECT 123.000 49.100 123.400 49.200 ;
        RECT 126.200 49.100 126.600 49.200 ;
        RECT 123.000 48.800 126.600 49.100 ;
        RECT 127.000 49.100 127.400 49.200 ;
        RECT 141.400 49.100 141.800 49.200 ;
        RECT 127.000 48.800 141.800 49.100 ;
        RECT 147.800 49.100 148.200 49.200 ;
        RECT 150.200 49.100 150.600 49.200 ;
        RECT 147.800 48.800 150.600 49.100 ;
        RECT 111.800 48.200 112.100 48.800 ;
        RECT 126.200 48.200 126.500 48.800 ;
        RECT 2.200 47.800 2.600 48.200 ;
        RECT 7.800 48.100 8.200 48.200 ;
        RECT 11.000 48.100 11.400 48.200 ;
        RECT 19.000 48.100 19.400 48.200 ;
        RECT 7.800 47.800 19.400 48.100 ;
        RECT 27.000 48.100 27.400 48.200 ;
        RECT 35.800 48.100 36.200 48.200 ;
        RECT 27.000 47.800 36.200 48.100 ;
        RECT 38.200 48.100 38.600 48.200 ;
        RECT 40.600 48.100 41.000 48.200 ;
        RECT 43.800 48.100 44.200 48.200 ;
        RECT 46.200 48.100 46.600 48.200 ;
        RECT 38.200 47.800 46.600 48.100 ;
        RECT 49.400 48.100 49.800 48.200 ;
        RECT 50.200 48.100 50.600 48.200 ;
        RECT 49.400 47.800 50.600 48.100 ;
        RECT 51.000 48.100 51.400 48.200 ;
        RECT 65.400 48.100 65.800 48.200 ;
        RECT 69.400 48.100 69.800 48.200 ;
        RECT 51.000 47.800 69.800 48.100 ;
        RECT 71.000 48.100 71.400 48.200 ;
        RECT 72.600 48.100 73.000 48.200 ;
        RECT 71.000 47.800 73.000 48.100 ;
        RECT 75.000 48.100 75.400 48.200 ;
        RECT 86.200 48.100 86.600 48.200 ;
        RECT 75.000 47.800 86.600 48.100 ;
        RECT 87.800 48.100 88.200 48.200 ;
        RECT 91.000 48.100 91.400 48.200 ;
        RECT 87.800 47.800 91.400 48.100 ;
        RECT 92.600 48.100 93.000 48.200 ;
        RECT 103.000 48.100 103.400 48.200 ;
        RECT 103.800 48.100 104.200 48.200 ;
        RECT 107.800 48.100 108.200 48.200 ;
        RECT 92.600 47.800 104.200 48.100 ;
        RECT 104.600 47.800 108.200 48.100 ;
        RECT 111.800 47.800 112.200 48.200 ;
        RECT 126.200 47.800 126.600 48.200 ;
        RECT 128.600 48.100 129.000 48.200 ;
        RECT 134.200 48.100 134.600 48.200 ;
        RECT 128.600 47.800 134.600 48.100 ;
        RECT 139.800 48.100 140.200 48.200 ;
        RECT 147.800 48.100 148.200 48.200 ;
        RECT 149.400 48.100 149.800 48.200 ;
        RECT 139.800 47.800 149.800 48.100 ;
        RECT 2.200 47.100 2.500 47.800 ;
        RECT 3.800 47.100 4.200 47.200 ;
        RECT 2.200 46.800 4.200 47.100 ;
        RECT 8.600 46.800 9.000 47.200 ;
        RECT 14.200 47.100 14.600 47.200 ;
        RECT 16.600 47.100 17.000 47.200 ;
        RECT 14.200 46.800 17.000 47.100 ;
        RECT 31.000 47.100 31.400 47.200 ;
        RECT 43.800 47.100 44.200 47.200 ;
        RECT 31.000 46.800 44.200 47.100 ;
        RECT 44.600 47.100 45.000 47.200 ;
        RECT 48.600 47.100 49.000 47.200 ;
        RECT 44.600 46.800 49.000 47.100 ;
        RECT 54.200 47.100 54.600 47.200 ;
        RECT 58.200 47.100 58.600 47.200 ;
        RECT 54.200 46.800 58.600 47.100 ;
        RECT 59.000 47.100 59.400 47.200 ;
        RECT 61.400 47.100 61.800 47.200 ;
        RECT 63.800 47.100 64.200 47.200 ;
        RECT 59.000 46.800 64.200 47.100 ;
        RECT 69.400 47.100 69.800 47.200 ;
        RECT 71.000 47.100 71.400 47.200 ;
        RECT 69.400 46.800 71.400 47.100 ;
        RECT 79.000 46.800 79.400 47.200 ;
        RECT 79.800 47.100 80.200 47.200 ;
        RECT 81.400 47.100 81.800 47.200 ;
        RECT 79.800 46.800 81.800 47.100 ;
        RECT 88.600 47.100 89.000 47.200 ;
        RECT 89.400 47.100 89.800 47.200 ;
        RECT 88.600 46.800 89.800 47.100 ;
        RECT 92.600 47.100 93.000 47.200 ;
        RECT 99.000 47.100 99.400 47.200 ;
        RECT 92.600 46.800 99.400 47.100 ;
        RECT 99.800 47.100 100.200 47.200 ;
        RECT 100.600 47.100 101.000 47.200 ;
        RECT 99.800 46.800 101.000 47.100 ;
        RECT 101.400 47.100 101.800 47.200 ;
        RECT 104.600 47.100 104.900 47.800 ;
        RECT 101.400 46.800 104.900 47.100 ;
        RECT 105.400 47.100 105.800 47.200 ;
        RECT 106.200 47.100 106.600 47.200 ;
        RECT 105.400 46.800 106.600 47.100 ;
        RECT 108.600 47.100 109.000 47.200 ;
        RECT 110.200 47.100 110.600 47.200 ;
        RECT 108.600 46.800 110.600 47.100 ;
        RECT 115.000 47.100 115.400 47.200 ;
        RECT 117.400 47.100 117.800 47.200 ;
        RECT 115.000 46.800 117.800 47.100 ;
        RECT 121.400 47.100 121.800 47.200 ;
        RECT 131.800 47.100 132.200 47.200 ;
        RECT 121.400 46.800 132.200 47.100 ;
        RECT 134.200 47.100 134.600 47.200 ;
        RECT 135.000 47.100 135.400 47.200 ;
        RECT 135.800 47.100 136.200 47.200 ;
        RECT 134.200 46.800 136.200 47.100 ;
        RECT 136.600 46.800 137.000 47.200 ;
        RECT 8.600 46.200 8.900 46.800 ;
        RECT 39.800 46.200 40.100 46.800 ;
        RECT 79.000 46.200 79.300 46.800 ;
        RECT 136.600 46.200 136.900 46.800 ;
        RECT 5.400 46.100 5.800 46.200 ;
        RECT 7.000 46.100 7.400 46.200 ;
        RECT 5.400 45.800 7.400 46.100 ;
        RECT 8.600 45.800 9.000 46.200 ;
        RECT 17.400 46.100 17.800 46.200 ;
        RECT 19.000 46.100 19.400 46.200 ;
        RECT 17.400 45.800 19.400 46.100 ;
        RECT 30.200 46.100 30.600 46.200 ;
        RECT 38.200 46.100 38.600 46.200 ;
        RECT 39.000 46.100 39.400 46.200 ;
        RECT 30.200 45.800 39.400 46.100 ;
        RECT 39.800 45.800 40.200 46.200 ;
        RECT 45.400 46.100 45.800 46.200 ;
        RECT 46.200 46.100 46.600 46.200 ;
        RECT 45.400 45.800 46.600 46.100 ;
        RECT 47.800 46.100 48.200 46.200 ;
        RECT 51.000 46.100 51.400 46.200 ;
        RECT 47.800 45.800 51.400 46.100 ;
        RECT 75.800 46.100 76.200 46.200 ;
        RECT 76.600 46.100 77.000 46.200 ;
        RECT 75.800 45.800 77.000 46.100 ;
        RECT 79.000 45.800 79.400 46.200 ;
        RECT 80.600 46.100 81.000 46.200 ;
        RECT 86.200 46.100 86.600 46.200 ;
        RECT 80.600 45.800 86.600 46.100 ;
        RECT 91.800 46.100 92.200 46.200 ;
        RECT 95.000 46.100 95.400 46.200 ;
        RECT 91.800 45.800 95.400 46.100 ;
        RECT 97.400 46.100 97.800 46.200 ;
        RECT 99.000 46.100 99.400 46.200 ;
        RECT 102.200 46.100 102.600 46.200 ;
        RECT 122.200 46.100 122.600 46.200 ;
        RECT 124.600 46.100 125.000 46.200 ;
        RECT 97.400 45.800 116.100 46.100 ;
        RECT 122.200 45.800 125.000 46.100 ;
        RECT 127.800 46.100 128.200 46.200 ;
        RECT 128.600 46.100 129.000 46.200 ;
        RECT 127.800 45.800 129.000 46.100 ;
        RECT 130.200 45.800 130.600 46.200 ;
        RECT 136.600 46.100 137.000 46.200 ;
        RECT 145.400 46.100 145.800 46.200 ;
        RECT 136.600 45.800 145.800 46.100 ;
        RECT 115.800 45.200 116.100 45.800 ;
        RECT 3.000 45.100 3.400 45.200 ;
        RECT 6.200 45.100 6.600 45.200 ;
        RECT 34.200 45.100 34.600 45.200 ;
        RECT 40.600 45.100 41.000 45.200 ;
        RECT 3.000 44.800 14.500 45.100 ;
        RECT 34.200 44.800 41.000 45.100 ;
        RECT 52.600 45.100 53.000 45.200 ;
        RECT 55.800 45.100 56.200 45.200 ;
        RECT 52.600 44.800 56.200 45.100 ;
        RECT 75.800 45.100 76.200 45.200 ;
        RECT 78.200 45.100 78.600 45.200 ;
        RECT 75.800 44.800 78.600 45.100 ;
        RECT 85.400 45.100 85.800 45.200 ;
        RECT 94.200 45.100 94.600 45.200 ;
        RECT 95.800 45.100 96.200 45.200 ;
        RECT 85.400 44.800 96.200 45.100 ;
        RECT 99.800 45.100 100.200 45.200 ;
        RECT 101.400 45.100 101.800 45.200 ;
        RECT 99.800 44.800 101.800 45.100 ;
        RECT 105.400 45.100 105.800 45.200 ;
        RECT 107.800 45.100 108.200 45.200 ;
        RECT 108.600 45.100 109.000 45.200 ;
        RECT 105.400 44.800 109.000 45.100 ;
        RECT 115.800 44.800 116.200 45.200 ;
        RECT 123.000 45.100 123.400 45.200 ;
        RECT 130.200 45.100 130.500 45.800 ;
        RECT 123.000 44.800 130.500 45.100 ;
        RECT 136.600 45.100 137.000 45.200 ;
        RECT 139.800 45.100 140.200 45.200 ;
        RECT 136.600 44.800 140.200 45.100 ;
        RECT 14.200 44.200 14.500 44.800 ;
        RECT 10.200 44.100 10.600 44.200 ;
        RECT 11.000 44.100 11.400 44.200 ;
        RECT 10.200 43.800 11.400 44.100 ;
        RECT 14.200 43.800 14.600 44.200 ;
        RECT 27.800 44.100 28.200 44.200 ;
        RECT 31.000 44.100 31.400 44.200 ;
        RECT 27.800 43.800 31.400 44.100 ;
        RECT 42.200 44.100 42.600 44.200 ;
        RECT 50.200 44.100 50.600 44.200 ;
        RECT 42.200 43.800 50.600 44.100 ;
        RECT 68.600 44.100 69.000 44.200 ;
        RECT 71.800 44.100 72.200 44.200 ;
        RECT 68.600 43.800 72.200 44.100 ;
        RECT 81.400 44.100 81.800 44.200 ;
        RECT 106.200 44.100 106.600 44.200 ;
        RECT 123.000 44.100 123.400 44.200 ;
        RECT 81.400 43.800 123.400 44.100 ;
        RECT 11.800 43.100 12.200 43.200 ;
        RECT 14.200 43.100 14.600 43.200 ;
        RECT 11.800 42.800 14.600 43.100 ;
        RECT 34.200 43.100 34.600 43.200 ;
        RECT 52.600 43.100 53.000 43.200 ;
        RECT 34.200 42.800 53.000 43.100 ;
        RECT 55.000 43.100 55.400 43.200 ;
        RECT 81.400 43.100 81.800 43.200 ;
        RECT 55.000 42.800 81.800 43.100 ;
        RECT 85.400 43.100 85.800 43.200 ;
        RECT 87.000 43.100 87.400 43.200 ;
        RECT 85.400 42.800 87.400 43.100 ;
        RECT 96.600 43.100 97.000 43.200 ;
        RECT 104.600 43.100 105.000 43.200 ;
        RECT 96.600 42.800 105.000 43.100 ;
        RECT 117.400 43.100 117.800 43.200 ;
        RECT 131.000 43.100 131.400 43.200 ;
        RECT 141.400 43.100 141.800 43.200 ;
        RECT 117.400 42.800 141.800 43.100 ;
        RECT 8.600 42.100 9.000 42.200 ;
        RECT 20.600 42.100 21.000 42.200 ;
        RECT 8.600 41.800 21.000 42.100 ;
        RECT 41.400 42.100 41.800 42.200 ;
        RECT 75.800 42.100 76.200 42.200 ;
        RECT 77.400 42.100 77.800 42.200 ;
        RECT 88.600 42.100 89.000 42.200 ;
        RECT 138.200 42.100 138.600 42.200 ;
        RECT 41.400 41.800 138.600 42.100 ;
        RECT 50.200 41.100 50.600 41.200 ;
        RECT 58.200 41.100 58.600 41.200 ;
        RECT 62.200 41.100 62.600 41.200 ;
        RECT 77.400 41.100 77.800 41.200 ;
        RECT 123.800 41.100 124.200 41.200 ;
        RECT 50.200 40.800 77.800 41.100 ;
        RECT 107.800 40.800 124.200 41.100 ;
        RECT 125.400 41.100 125.800 41.200 ;
        RECT 127.000 41.100 127.400 41.200 ;
        RECT 133.400 41.100 133.800 41.200 ;
        RECT 135.800 41.100 136.200 41.200 ;
        RECT 125.400 40.800 136.200 41.100 ;
        RECT 136.600 41.100 137.000 41.200 ;
        RECT 140.600 41.100 141.000 41.200 ;
        RECT 136.600 40.800 141.000 41.100 ;
        RECT 51.800 40.100 52.200 40.200 ;
        RECT 59.800 40.100 60.200 40.200 ;
        RECT 51.800 39.800 60.200 40.100 ;
        RECT 61.400 40.100 61.800 40.200 ;
        RECT 69.400 40.100 69.800 40.200 ;
        RECT 61.400 39.800 69.800 40.100 ;
        RECT 76.600 40.100 77.000 40.200 ;
        RECT 107.800 40.100 108.100 40.800 ;
        RECT 76.600 39.800 108.100 40.100 ;
        RECT 108.600 40.100 109.000 40.200 ;
        RECT 113.400 40.100 113.800 40.200 ;
        RECT 108.600 39.800 113.800 40.100 ;
        RECT 115.800 40.100 116.200 40.200 ;
        RECT 121.400 40.100 121.800 40.200 ;
        RECT 115.800 39.800 121.800 40.100 ;
        RECT 132.600 40.100 133.000 40.200 ;
        RECT 133.400 40.100 133.800 40.200 ;
        RECT 132.600 39.800 133.800 40.100 ;
        RECT 19.000 39.100 19.400 39.200 ;
        RECT 27.800 39.100 28.200 39.200 ;
        RECT 55.000 39.100 55.400 39.200 ;
        RECT 19.000 38.800 28.200 39.100 ;
        RECT 39.800 38.800 55.400 39.100 ;
        RECT 55.800 39.100 56.200 39.200 ;
        RECT 71.800 39.100 72.200 39.200 ;
        RECT 79.800 39.100 80.200 39.200 ;
        RECT 86.200 39.100 86.600 39.200 ;
        RECT 91.800 39.100 92.200 39.200 ;
        RECT 112.600 39.100 113.000 39.200 ;
        RECT 55.800 38.800 113.000 39.100 ;
        RECT 119.800 39.100 120.200 39.200 ;
        RECT 119.800 38.800 128.900 39.100 ;
        RECT 39.800 38.200 40.100 38.800 ;
        RECT 128.600 38.200 128.900 38.800 ;
        RECT 15.000 38.100 15.400 38.200 ;
        RECT 21.400 38.100 21.800 38.200 ;
        RECT 15.000 37.800 21.800 38.100 ;
        RECT 39.800 37.800 40.200 38.200 ;
        RECT 59.000 38.100 59.400 38.200 ;
        RECT 57.400 37.800 59.400 38.100 ;
        RECT 60.600 38.100 61.000 38.200 ;
        RECT 84.600 38.100 85.000 38.200 ;
        RECT 60.600 37.800 85.000 38.100 ;
        RECT 94.200 38.100 94.600 38.200 ;
        RECT 104.600 38.100 105.000 38.200 ;
        RECT 107.000 38.100 107.400 38.200 ;
        RECT 94.200 37.800 107.400 38.100 ;
        RECT 107.800 38.100 108.200 38.200 ;
        RECT 110.200 38.100 110.600 38.200 ;
        RECT 107.800 37.800 110.600 38.100 ;
        RECT 128.600 37.800 129.000 38.200 ;
        RECT 57.400 37.200 57.700 37.800 ;
        RECT 7.800 36.800 8.200 37.200 ;
        RECT 12.600 36.800 13.000 37.200 ;
        RECT 18.200 37.100 18.600 37.200 ;
        RECT 20.600 37.100 21.000 37.200 ;
        RECT 18.200 36.800 21.000 37.100 ;
        RECT 35.000 37.100 35.400 37.200 ;
        RECT 41.400 37.100 41.800 37.200 ;
        RECT 35.000 36.800 41.800 37.100 ;
        RECT 57.400 36.800 57.800 37.200 ;
        RECT 59.800 37.100 60.200 37.200 ;
        RECT 80.600 37.100 81.000 37.200 ;
        RECT 83.800 37.100 84.200 37.200 ;
        RECT 59.800 36.800 84.200 37.100 ;
        RECT 87.800 37.100 88.200 37.200 ;
        RECT 95.800 37.100 96.200 37.200 ;
        RECT 87.800 36.800 96.200 37.100 ;
        RECT 101.400 37.100 101.800 37.200 ;
        RECT 106.200 37.100 106.600 37.200 ;
        RECT 117.400 37.100 117.800 37.200 ;
        RECT 101.400 36.800 117.800 37.100 ;
        RECT 7.800 36.200 8.100 36.800 ;
        RECT 7.800 35.800 8.200 36.200 ;
        RECT 8.600 35.800 9.000 36.200 ;
        RECT 12.600 36.100 12.900 36.800 ;
        RECT 25.400 36.100 25.800 36.200 ;
        RECT 12.600 35.800 25.800 36.100 ;
        RECT 73.400 36.100 73.800 36.200 ;
        RECT 82.200 36.100 82.600 36.200 ;
        RECT 73.400 35.800 82.600 36.100 ;
        RECT 83.800 36.100 84.200 36.200 ;
        RECT 87.000 36.100 87.400 36.200 ;
        RECT 83.800 35.800 87.400 36.100 ;
        RECT 90.200 36.100 90.600 36.200 ;
        RECT 92.600 36.100 93.000 36.200 ;
        RECT 90.200 35.800 93.000 36.100 ;
        RECT 104.600 36.100 105.000 36.200 ;
        RECT 107.800 36.100 108.200 36.200 ;
        RECT 104.600 35.800 108.200 36.100 ;
        RECT 108.600 36.100 109.000 36.200 ;
        RECT 111.000 36.100 111.400 36.200 ;
        RECT 108.600 35.800 111.400 36.100 ;
        RECT 138.200 36.100 138.600 36.200 ;
        RECT 139.000 36.100 139.400 36.200 ;
        RECT 143.800 36.100 144.200 36.200 ;
        RECT 138.200 35.800 144.200 36.100 ;
        RECT 8.600 35.200 8.900 35.800 ;
        RECT 2.200 35.100 2.600 35.200 ;
        RECT 3.000 35.100 3.400 35.200 ;
        RECT 2.200 34.800 3.400 35.100 ;
        RECT 4.600 35.100 5.000 35.200 ;
        RECT 7.000 35.100 7.400 35.200 ;
        RECT 4.600 34.800 7.400 35.100 ;
        RECT 8.600 34.800 9.000 35.200 ;
        RECT 10.200 35.100 10.600 35.200 ;
        RECT 16.600 35.100 17.000 35.200 ;
        RECT 10.200 34.800 17.000 35.100 ;
        RECT 21.400 35.100 21.800 35.200 ;
        RECT 23.000 35.100 23.400 35.200 ;
        RECT 21.400 34.800 23.400 35.100 ;
        RECT 37.400 35.100 37.800 35.200 ;
        RECT 47.800 35.100 48.200 35.200 ;
        RECT 64.600 35.100 65.000 35.200 ;
        RECT 37.400 34.800 65.000 35.100 ;
        RECT 70.200 35.100 70.600 35.200 ;
        RECT 71.000 35.100 71.400 35.200 ;
        RECT 70.200 34.800 71.400 35.100 ;
        RECT 73.400 35.100 73.800 35.200 ;
        RECT 75.000 35.100 75.400 35.200 ;
        RECT 73.400 34.800 75.400 35.100 ;
        RECT 81.400 34.800 81.800 35.200 ;
        RECT 83.000 35.100 83.400 35.200 ;
        RECT 82.200 34.800 83.400 35.100 ;
        RECT 83.800 35.100 84.200 35.200 ;
        RECT 84.600 35.100 85.000 35.200 ;
        RECT 83.800 34.800 85.000 35.100 ;
        RECT 86.200 35.100 86.600 35.200 ;
        RECT 91.000 35.100 91.400 35.200 ;
        RECT 103.000 35.100 103.400 35.200 ;
        RECT 86.200 34.800 103.400 35.100 ;
        RECT 104.600 35.100 105.000 35.200 ;
        RECT 109.400 35.100 109.800 35.200 ;
        RECT 104.600 34.800 109.800 35.100 ;
        RECT 111.800 35.100 112.200 35.200 ;
        RECT 115.000 35.100 115.400 35.200 ;
        RECT 111.800 34.800 115.400 35.100 ;
        RECT 119.800 35.100 120.200 35.200 ;
        RECT 123.800 35.100 124.200 35.200 ;
        RECT 119.800 34.800 124.200 35.100 ;
        RECT 134.200 35.100 134.600 35.200 ;
        RECT 135.800 35.100 136.200 35.200 ;
        RECT 137.400 35.100 137.800 35.200 ;
        RECT 134.200 34.800 137.800 35.100 ;
        RECT 140.600 35.100 141.000 35.200 ;
        RECT 143.000 35.100 143.400 35.200 ;
        RECT 140.600 34.800 143.400 35.100 ;
        RECT 81.400 34.200 81.700 34.800 ;
        RECT 82.200 34.200 82.500 34.800 ;
        RECT 3.800 34.100 4.200 34.200 ;
        RECT 6.200 34.100 6.600 34.200 ;
        RECT 7.800 34.100 8.200 34.200 ;
        RECT 15.000 34.100 15.400 34.200 ;
        RECT 3.800 33.800 5.700 34.100 ;
        RECT 6.200 33.800 8.200 34.100 ;
        RECT 10.200 33.800 15.400 34.100 ;
        RECT 15.800 34.100 16.200 34.200 ;
        RECT 36.600 34.100 37.000 34.200 ;
        RECT 15.800 33.800 37.000 34.100 ;
        RECT 69.400 34.100 69.800 34.200 ;
        RECT 79.800 34.100 80.200 34.200 ;
        RECT 69.400 33.800 80.200 34.100 ;
        RECT 81.400 33.800 81.800 34.200 ;
        RECT 82.200 33.800 82.600 34.200 ;
        RECT 83.000 34.100 83.400 34.200 ;
        RECT 88.600 34.100 89.000 34.200 ;
        RECT 91.800 34.100 92.200 34.200 ;
        RECT 126.200 34.100 126.600 34.200 ;
        RECT 83.000 33.800 126.600 34.100 ;
        RECT 140.600 34.100 141.000 34.200 ;
        RECT 142.200 34.100 142.600 34.200 ;
        RECT 147.800 34.100 148.200 34.200 ;
        RECT 140.600 33.800 148.200 34.100 ;
        RECT 5.400 33.200 5.700 33.800 ;
        RECT 10.200 33.200 10.500 33.800 ;
        RECT 5.400 32.800 5.800 33.200 ;
        RECT 10.200 32.800 10.600 33.200 ;
        RECT 17.400 33.100 17.800 33.200 ;
        RECT 20.600 33.100 21.000 33.200 ;
        RECT 17.400 32.800 21.000 33.100 ;
        RECT 32.600 33.100 33.000 33.200 ;
        RECT 36.600 33.100 37.000 33.200 ;
        RECT 32.600 32.800 37.000 33.100 ;
        RECT 65.400 33.100 65.800 33.200 ;
        RECT 71.800 33.100 72.200 33.200 ;
        RECT 65.400 32.800 72.200 33.100 ;
        RECT 74.200 32.800 74.600 33.200 ;
        RECT 75.000 32.800 75.400 33.200 ;
        RECT 84.600 33.100 85.000 33.200 ;
        RECT 88.600 33.100 89.000 33.200 ;
        RECT 83.800 32.800 89.000 33.100 ;
        RECT 111.000 33.100 111.400 33.200 ;
        RECT 111.800 33.100 112.200 33.200 ;
        RECT 111.000 32.800 112.200 33.100 ;
        RECT 118.200 32.800 118.600 33.200 ;
        RECT 128.600 33.100 129.000 33.200 ;
        RECT 129.400 33.100 129.800 33.200 ;
        RECT 128.600 32.800 129.800 33.100 ;
        RECT 133.400 33.100 133.800 33.200 ;
        RECT 138.200 33.100 138.600 33.200 ;
        RECT 133.400 32.800 138.600 33.100 ;
        RECT 74.200 32.200 74.500 32.800 ;
        RECT 75.000 32.200 75.300 32.800 ;
        RECT 7.000 32.100 7.400 32.200 ;
        RECT 13.400 32.100 13.800 32.200 ;
        RECT 7.000 31.800 13.800 32.100 ;
        RECT 14.200 32.100 14.600 32.200 ;
        RECT 19.000 32.100 19.400 32.200 ;
        RECT 14.200 31.800 19.400 32.100 ;
        RECT 74.200 31.800 74.600 32.200 ;
        RECT 75.000 31.800 75.400 32.200 ;
        RECT 87.800 32.100 88.200 32.200 ;
        RECT 98.200 32.100 98.600 32.200 ;
        RECT 87.800 31.800 98.600 32.100 ;
        RECT 109.400 32.100 109.800 32.200 ;
        RECT 111.000 32.100 111.400 32.200 ;
        RECT 109.400 31.800 111.400 32.100 ;
        RECT 118.200 32.100 118.500 32.800 ;
        RECT 131.800 32.100 132.200 32.200 ;
        RECT 118.200 31.800 132.200 32.100 ;
        RECT 4.600 31.100 5.000 31.200 ;
        RECT 7.800 31.100 8.200 31.200 ;
        RECT 10.200 31.100 10.600 31.200 ;
        RECT 4.600 30.800 10.600 31.100 ;
        RECT 75.000 31.100 75.400 31.200 ;
        RECT 78.200 31.100 78.600 31.200 ;
        RECT 84.600 31.100 85.000 31.200 ;
        RECT 75.000 30.800 85.000 31.100 ;
        RECT 109.400 31.100 109.800 31.200 ;
        RECT 120.600 31.100 121.000 31.200 ;
        RECT 121.400 31.100 121.800 31.200 ;
        RECT 109.400 30.800 121.800 31.100 ;
        RECT 23.800 30.100 24.200 30.200 ;
        RECT 28.600 30.100 29.000 30.200 ;
        RECT 23.800 29.800 29.000 30.100 ;
        RECT 44.600 30.100 45.000 30.200 ;
        RECT 60.600 30.100 61.000 30.200 ;
        RECT 62.200 30.100 62.600 30.200 ;
        RECT 44.600 29.800 62.600 30.100 ;
        RECT 64.600 30.100 65.000 30.200 ;
        RECT 81.400 30.100 81.800 30.200 ;
        RECT 87.000 30.100 87.400 30.200 ;
        RECT 64.600 29.800 87.400 30.100 ;
        RECT 95.800 30.100 96.200 30.200 ;
        RECT 99.000 30.100 99.400 30.200 ;
        RECT 95.800 29.800 99.400 30.100 ;
        RECT 103.800 30.100 104.200 30.200 ;
        RECT 112.600 30.100 113.000 30.200 ;
        RECT 103.800 29.800 113.000 30.100 ;
        RECT 119.000 30.100 119.400 30.200 ;
        RECT 122.200 30.100 122.600 30.200 ;
        RECT 128.600 30.100 129.000 30.200 ;
        RECT 119.000 29.800 129.000 30.100 ;
        RECT 0.600 29.100 1.000 29.200 ;
        RECT 15.800 29.100 16.200 29.200 ;
        RECT 0.600 28.800 16.200 29.100 ;
        RECT 38.200 29.100 38.600 29.200 ;
        RECT 40.600 29.100 41.000 29.200 ;
        RECT 45.400 29.100 45.800 29.200 ;
        RECT 46.200 29.100 46.600 29.200 ;
        RECT 38.200 28.800 46.600 29.100 ;
        RECT 59.000 29.100 59.400 29.200 ;
        RECT 65.400 29.100 65.800 29.200 ;
        RECT 69.400 29.100 69.800 29.200 ;
        RECT 59.000 28.800 69.800 29.100 ;
        RECT 73.400 29.100 73.800 29.200 ;
        RECT 77.400 29.100 77.800 29.200 ;
        RECT 73.400 28.800 77.800 29.100 ;
        RECT 78.200 28.800 78.600 29.200 ;
        RECT 79.000 29.100 79.400 29.200 ;
        RECT 85.400 29.100 85.800 29.200 ;
        RECT 109.400 29.100 109.800 29.200 ;
        RECT 79.000 28.800 85.800 29.100 ;
        RECT 86.200 28.800 109.800 29.100 ;
        RECT 114.200 28.800 114.600 29.200 ;
        RECT 115.000 29.100 115.400 29.200 ;
        RECT 117.400 29.100 117.800 29.200 ;
        RECT 115.000 28.800 117.800 29.100 ;
        RECT 121.400 29.100 121.800 29.200 ;
        RECT 125.400 29.100 125.800 29.200 ;
        RECT 121.400 28.800 125.800 29.100 ;
        RECT 126.200 29.100 126.600 29.200 ;
        RECT 139.800 29.100 140.200 29.200 ;
        RECT 126.200 28.800 140.200 29.100 ;
        RECT 5.400 28.100 5.800 28.200 ;
        RECT 9.400 28.100 9.800 28.200 ;
        RECT 5.400 27.800 9.800 28.100 ;
        RECT 39.000 28.100 39.400 28.200 ;
        RECT 50.200 28.100 50.600 28.200 ;
        RECT 39.000 27.800 50.600 28.100 ;
        RECT 62.200 28.100 62.600 28.200 ;
        RECT 67.800 28.100 68.200 28.200 ;
        RECT 62.200 27.800 68.200 28.100 ;
        RECT 68.600 28.100 69.000 28.200 ;
        RECT 70.200 28.100 70.600 28.200 ;
        RECT 68.600 27.800 70.600 28.100 ;
        RECT 71.000 28.100 71.400 28.200 ;
        RECT 78.200 28.100 78.500 28.800 ;
        RECT 86.200 28.200 86.500 28.800 ;
        RECT 80.600 28.100 81.000 28.200 ;
        RECT 83.800 28.100 84.200 28.200 ;
        RECT 71.000 27.800 76.900 28.100 ;
        RECT 78.200 27.800 84.200 28.100 ;
        RECT 86.200 27.800 86.600 28.200 ;
        RECT 91.800 28.100 92.200 28.200 ;
        RECT 95.800 28.100 96.200 28.200 ;
        RECT 91.800 27.800 96.200 28.100 ;
        RECT 97.400 28.100 97.800 28.200 ;
        RECT 109.400 28.100 109.800 28.200 ;
        RECT 97.400 27.800 109.800 28.100 ;
        RECT 110.200 28.100 110.600 28.200 ;
        RECT 114.200 28.100 114.500 28.800 ;
        RECT 110.200 27.800 114.500 28.100 ;
        RECT 115.800 28.100 116.200 28.200 ;
        RECT 127.000 28.100 127.400 28.200 ;
        RECT 115.800 27.800 127.400 28.100 ;
        RECT 13.400 27.100 13.800 27.200 ;
        RECT 17.400 27.100 17.800 27.200 ;
        RECT 13.400 26.800 17.800 27.100 ;
        RECT 21.400 27.100 21.800 27.200 ;
        RECT 27.000 27.100 27.400 27.200 ;
        RECT 21.400 26.800 27.400 27.100 ;
        RECT 30.200 27.100 30.600 27.200 ;
        RECT 41.400 27.100 41.800 27.200 ;
        RECT 47.000 27.100 47.400 27.200 ;
        RECT 30.200 26.800 47.400 27.100 ;
        RECT 56.600 26.800 57.000 27.200 ;
        RECT 61.400 27.100 61.800 27.200 ;
        RECT 73.400 27.100 73.800 27.200 ;
        RECT 61.400 26.800 73.800 27.100 ;
        RECT 75.800 26.800 76.200 27.200 ;
        RECT 76.600 27.100 76.900 27.800 ;
        RECT 89.400 27.100 89.800 27.200 ;
        RECT 91.000 27.100 91.400 27.200 ;
        RECT 76.600 26.800 91.400 27.100 ;
        RECT 92.600 26.800 93.000 27.200 ;
        RECT 94.200 27.100 94.600 27.200 ;
        RECT 95.000 27.100 95.400 27.200 ;
        RECT 94.200 26.800 95.400 27.100 ;
        RECT 97.400 27.100 97.800 27.200 ;
        RECT 98.200 27.100 98.600 27.200 ;
        RECT 97.400 26.800 98.600 27.100 ;
        RECT 100.600 27.100 101.000 27.200 ;
        RECT 105.400 27.100 105.800 27.200 ;
        RECT 106.200 27.100 106.600 27.200 ;
        RECT 100.600 27.000 103.300 27.100 ;
        RECT 100.600 26.800 103.400 27.000 ;
        RECT 105.400 26.800 106.600 27.100 ;
        RECT 107.800 27.100 108.200 27.200 ;
        RECT 108.600 27.100 109.000 27.200 ;
        RECT 107.800 26.800 109.000 27.100 ;
        RECT 111.800 27.100 112.200 27.200 ;
        RECT 112.600 27.100 113.000 27.200 ;
        RECT 111.800 26.800 113.000 27.100 ;
        RECT 115.000 27.100 115.400 27.200 ;
        RECT 115.800 27.100 116.200 27.200 ;
        RECT 115.000 26.800 116.200 27.100 ;
        RECT 116.600 27.100 117.000 27.200 ;
        RECT 119.000 27.100 119.400 27.200 ;
        RECT 116.600 26.800 119.400 27.100 ;
        RECT 123.000 27.100 123.400 27.200 ;
        RECT 123.800 27.100 124.200 27.200 ;
        RECT 123.000 26.800 124.200 27.100 ;
        RECT 125.400 27.100 125.800 27.200 ;
        RECT 129.400 27.100 129.800 27.200 ;
        RECT 136.600 27.100 137.000 27.200 ;
        RECT 125.400 26.800 127.300 27.100 ;
        RECT 129.400 26.800 137.000 27.100 ;
        RECT 142.200 27.100 142.600 27.200 ;
        RECT 145.400 27.100 145.800 27.200 ;
        RECT 142.200 26.800 145.800 27.100 ;
        RECT 2.200 26.100 2.600 26.200 ;
        RECT 7.000 26.100 7.400 26.200 ;
        RECT 8.600 26.100 9.000 26.200 ;
        RECT 18.200 26.100 18.600 26.200 ;
        RECT 19.800 26.100 20.200 26.200 ;
        RECT 2.200 25.800 9.000 26.100 ;
        RECT 16.600 25.800 20.200 26.100 ;
        RECT 42.200 26.100 42.600 26.200 ;
        RECT 44.600 26.100 45.000 26.200 ;
        RECT 46.200 26.100 46.600 26.200 ;
        RECT 42.200 25.800 46.600 26.100 ;
        RECT 56.600 26.100 56.900 26.800 ;
        RECT 75.800 26.200 76.100 26.800 ;
        RECT 57.400 26.100 57.800 26.200 ;
        RECT 56.600 25.800 57.800 26.100 ;
        RECT 59.000 25.800 59.400 26.200 ;
        RECT 67.000 26.100 67.400 26.200 ;
        RECT 71.000 26.100 71.400 26.200 ;
        RECT 67.000 25.800 71.400 26.100 ;
        RECT 75.800 25.800 76.200 26.200 ;
        RECT 76.600 25.800 77.000 26.200 ;
        RECT 92.600 26.100 92.900 26.800 ;
        RECT 103.000 26.600 103.400 26.800 ;
        RECT 127.000 26.200 127.300 26.800 ;
        RECT 99.000 26.100 99.400 26.200 ;
        RECT 116.600 26.100 117.000 26.200 ;
        RECT 92.600 25.800 117.000 26.100 ;
        RECT 124.600 26.100 125.000 26.200 ;
        RECT 126.200 26.100 126.600 26.200 ;
        RECT 124.600 25.800 126.600 26.100 ;
        RECT 127.000 26.100 127.400 26.200 ;
        RECT 130.200 26.100 130.600 26.200 ;
        RECT 133.400 26.100 133.800 26.200 ;
        RECT 127.000 25.800 133.800 26.100 ;
        RECT 139.000 26.100 139.400 26.200 ;
        RECT 141.400 26.100 141.800 26.200 ;
        RECT 139.000 25.800 141.800 26.100 ;
        RECT 16.600 25.200 16.900 25.800 ;
        RECT 3.800 25.100 4.200 25.200 ;
        RECT 7.800 25.100 8.200 25.200 ;
        RECT 11.800 25.100 12.200 25.200 ;
        RECT 3.800 24.800 12.200 25.100 ;
        RECT 16.600 24.800 17.000 25.200 ;
        RECT 55.800 25.100 56.200 25.200 ;
        RECT 59.000 25.100 59.300 25.800 ;
        RECT 76.600 25.200 76.900 25.800 ;
        RECT 63.000 25.100 63.400 25.200 ;
        RECT 34.200 24.800 43.300 25.100 ;
        RECT 55.800 24.800 63.400 25.100 ;
        RECT 68.600 25.100 69.000 25.200 ;
        RECT 75.000 25.100 75.400 25.200 ;
        RECT 75.800 25.100 76.200 25.200 ;
        RECT 68.600 24.800 76.200 25.100 ;
        RECT 76.600 24.800 77.000 25.200 ;
        RECT 85.400 25.100 85.800 25.200 ;
        RECT 107.000 25.100 107.400 25.200 ;
        RECT 109.400 25.100 109.800 25.200 ;
        RECT 85.400 24.800 109.800 25.100 ;
        RECT 117.400 25.100 117.800 25.200 ;
        RECT 119.800 25.100 120.200 25.200 ;
        RECT 117.400 24.800 120.200 25.100 ;
        RECT 122.200 25.100 122.600 25.200 ;
        RECT 146.200 25.100 146.600 25.200 ;
        RECT 122.200 24.800 146.600 25.100 ;
        RECT 34.200 24.200 34.500 24.800 ;
        RECT 43.000 24.200 43.300 24.800 ;
        RECT 8.600 24.100 9.000 24.200 ;
        RECT 10.200 24.100 10.600 24.200 ;
        RECT 8.600 23.800 10.600 24.100 ;
        RECT 15.800 24.100 16.200 24.200 ;
        RECT 19.800 24.100 20.200 24.200 ;
        RECT 25.400 24.100 25.800 24.200 ;
        RECT 15.800 23.800 25.800 24.100 ;
        RECT 34.200 23.800 34.600 24.200 ;
        RECT 43.000 24.100 43.400 24.200 ;
        RECT 53.400 24.100 53.800 24.200 ;
        RECT 54.200 24.100 54.600 24.200 ;
        RECT 43.000 23.800 54.600 24.100 ;
        RECT 65.400 24.100 65.800 24.200 ;
        RECT 82.200 24.100 82.600 24.200 ;
        RECT 65.400 23.800 82.600 24.100 ;
        RECT 92.600 24.100 93.000 24.200 ;
        RECT 93.400 24.100 93.800 24.200 ;
        RECT 92.600 23.800 93.800 24.100 ;
        RECT 104.600 24.100 105.000 24.200 ;
        RECT 113.400 24.100 113.800 24.200 ;
        RECT 104.600 23.800 113.800 24.100 ;
        RECT 51.000 23.100 51.400 23.200 ;
        RECT 58.200 23.100 58.600 23.200 ;
        RECT 51.000 22.800 58.600 23.100 ;
        RECT 80.600 23.100 81.000 23.200 ;
        RECT 94.200 23.100 94.600 23.200 ;
        RECT 80.600 22.800 94.600 23.100 ;
        RECT 107.000 23.100 107.400 23.200 ;
        RECT 122.200 23.100 122.600 23.200 ;
        RECT 139.000 23.100 139.400 23.200 ;
        RECT 143.000 23.100 143.400 23.200 ;
        RECT 107.000 22.800 143.400 23.100 ;
        RECT 35.000 22.100 35.400 22.200 ;
        RECT 37.400 22.100 37.800 22.200 ;
        RECT 35.000 21.800 37.800 22.100 ;
        RECT 56.600 22.100 57.000 22.200 ;
        RECT 74.200 22.100 74.600 22.200 ;
        RECT 80.600 22.100 81.000 22.200 ;
        RECT 56.600 21.800 81.000 22.100 ;
        RECT 88.600 22.100 89.000 22.200 ;
        RECT 103.800 22.100 104.200 22.200 ;
        RECT 88.600 21.800 104.200 22.100 ;
        RECT 112.600 22.100 113.000 22.200 ;
        RECT 126.200 22.100 126.600 22.200 ;
        RECT 112.600 21.800 126.600 22.100 ;
        RECT 79.800 21.100 80.200 21.200 ;
        RECT 107.800 21.100 108.200 21.200 ;
        RECT 111.800 21.100 112.200 21.200 ;
        RECT 124.600 21.100 125.000 21.200 ;
        RECT 79.800 20.800 125.000 21.100 ;
        RECT 126.200 21.100 126.600 21.200 ;
        RECT 128.600 21.100 129.000 21.200 ;
        RECT 126.200 20.800 129.000 21.100 ;
        RECT 77.400 20.100 77.800 20.200 ;
        RECT 103.800 20.100 104.200 20.200 ;
        RECT 108.600 20.100 109.000 20.200 ;
        RECT 77.400 19.800 109.000 20.100 ;
        RECT 113.400 20.100 113.800 20.200 ;
        RECT 123.000 20.100 123.400 20.200 ;
        RECT 113.400 19.800 123.400 20.100 ;
        RECT 133.400 19.800 133.800 20.200 ;
        RECT 18.200 19.100 18.600 19.200 ;
        RECT 18.200 18.800 20.100 19.100 ;
        RECT 19.800 18.200 20.100 18.800 ;
        RECT 74.200 18.800 74.600 19.200 ;
        RECT 108.600 19.100 108.900 19.800 ;
        RECT 133.400 19.200 133.700 19.800 ;
        RECT 127.000 19.100 127.400 19.200 ;
        RECT 132.600 19.100 133.000 19.200 ;
        RECT 108.600 18.800 133.000 19.100 ;
        RECT 133.400 18.800 133.800 19.200 ;
        RECT 1.400 18.100 1.800 18.200 ;
        RECT 1.400 17.800 15.300 18.100 ;
        RECT 19.800 17.800 20.200 18.200 ;
        RECT 24.600 18.100 25.000 18.200 ;
        RECT 31.000 18.100 31.400 18.200 ;
        RECT 32.600 18.100 33.000 18.200 ;
        RECT 24.600 17.800 33.000 18.100 ;
        RECT 34.200 17.800 34.600 18.200 ;
        RECT 72.600 18.100 73.000 18.200 ;
        RECT 74.200 18.100 74.500 18.800 ;
        RECT 72.600 17.800 74.500 18.100 ;
        RECT 94.200 18.100 94.600 18.200 ;
        RECT 95.800 18.100 96.200 18.200 ;
        RECT 94.200 17.800 96.200 18.100 ;
        RECT 98.200 18.100 98.600 18.200 ;
        RECT 114.200 18.100 114.600 18.200 ;
        RECT 121.400 18.100 121.800 18.200 ;
        RECT 134.200 18.100 134.600 18.200 ;
        RECT 140.600 18.100 141.000 18.200 ;
        RECT 98.200 17.800 141.000 18.100 ;
        RECT 15.000 17.200 15.300 17.800 ;
        RECT 6.200 16.800 6.600 17.200 ;
        RECT 15.000 16.800 15.400 17.200 ;
        RECT 16.600 17.100 17.000 17.200 ;
        RECT 34.200 17.100 34.500 17.800 ;
        RECT 16.600 16.800 34.500 17.100 ;
        RECT 36.600 17.100 37.000 17.200 ;
        RECT 39.800 17.100 40.200 17.200 ;
        RECT 36.600 16.800 40.200 17.100 ;
        RECT 44.600 17.100 45.000 17.200 ;
        RECT 53.400 17.100 53.800 17.200 ;
        RECT 44.600 16.800 53.800 17.100 ;
        RECT 55.800 16.800 56.200 17.200 ;
        RECT 75.000 17.100 75.400 17.200 ;
        RECT 92.600 17.100 93.000 17.200 ;
        RECT 75.000 16.800 93.000 17.100 ;
        RECT 95.800 17.100 96.200 17.200 ;
        RECT 106.200 17.100 106.600 17.200 ;
        RECT 95.800 16.800 106.600 17.100 ;
        RECT 115.000 17.100 115.400 17.200 ;
        RECT 126.200 17.100 126.600 17.200 ;
        RECT 115.000 16.800 126.600 17.100 ;
        RECT 127.800 17.100 128.200 17.200 ;
        RECT 128.600 17.100 129.000 17.200 ;
        RECT 135.800 17.100 136.200 17.200 ;
        RECT 127.800 16.800 136.200 17.100 ;
        RECT 2.200 15.800 2.600 16.200 ;
        RECT 3.800 15.800 4.200 16.200 ;
        RECT 6.200 16.100 6.500 16.800 ;
        RECT 10.200 16.100 10.600 16.200 ;
        RECT 6.200 15.800 10.600 16.100 ;
        RECT 14.200 16.100 14.600 16.200 ;
        RECT 16.600 16.100 17.000 16.200 ;
        RECT 14.200 15.800 17.000 16.100 ;
        RECT 18.200 16.100 18.600 16.200 ;
        RECT 21.400 16.100 21.800 16.200 ;
        RECT 18.200 15.800 21.800 16.100 ;
        RECT 27.800 16.100 28.200 16.200 ;
        RECT 31.800 16.100 32.200 16.200 ;
        RECT 27.800 15.800 32.200 16.100 ;
        RECT 35.000 15.800 35.400 16.200 ;
        RECT 36.600 16.100 37.000 16.200 ;
        RECT 40.600 16.100 41.000 16.200 ;
        RECT 43.800 16.100 44.200 16.200 ;
        RECT 36.600 15.800 44.200 16.100 ;
        RECT 45.400 16.100 45.800 16.200 ;
        RECT 48.600 16.100 49.000 16.200 ;
        RECT 55.800 16.100 56.100 16.800 ;
        RECT 45.400 15.800 56.100 16.100 ;
        RECT 63.800 16.100 64.200 16.200 ;
        RECT 67.800 16.100 68.200 16.200 ;
        RECT 63.800 15.800 68.200 16.100 ;
        RECT 75.000 16.100 75.400 16.200 ;
        RECT 76.600 16.100 77.000 16.200 ;
        RECT 75.000 15.800 77.000 16.100 ;
        RECT 77.400 16.100 77.800 16.200 ;
        RECT 85.400 16.100 85.800 16.200 ;
        RECT 77.400 15.800 85.800 16.100 ;
        RECT 87.800 16.100 88.200 16.200 ;
        RECT 106.200 16.100 106.600 16.200 ;
        RECT 87.800 15.800 106.600 16.100 ;
        RECT 107.000 16.100 107.400 16.200 ;
        RECT 108.600 16.100 109.000 16.200 ;
        RECT 107.000 15.800 109.000 16.100 ;
        RECT 110.200 16.100 110.600 16.200 ;
        RECT 113.400 16.100 113.800 16.200 ;
        RECT 110.200 15.800 113.800 16.100 ;
        RECT 121.400 16.100 121.800 16.200 ;
        RECT 122.200 16.100 122.600 16.200 ;
        RECT 121.400 15.800 122.600 16.100 ;
        RECT 136.600 16.100 137.000 16.200 ;
        RECT 139.000 16.100 139.400 16.200 ;
        RECT 136.600 15.800 139.400 16.100 ;
        RECT 147.800 16.100 148.200 16.200 ;
        RECT 148.600 16.100 149.000 16.200 ;
        RECT 147.800 15.800 149.000 16.100 ;
        RECT 2.200 15.100 2.500 15.800 ;
        RECT 3.800 15.100 4.100 15.800 ;
        RECT 2.200 14.800 4.100 15.100 ;
        RECT 6.200 15.100 6.600 15.200 ;
        RECT 13.400 15.100 13.800 15.200 ;
        RECT 23.000 15.100 23.400 15.200 ;
        RECT 29.400 15.100 29.800 15.200 ;
        RECT 35.000 15.100 35.300 15.800 ;
        RECT 6.200 14.800 35.300 15.100 ;
        RECT 66.200 15.100 66.600 15.200 ;
        RECT 70.200 15.100 70.600 15.200 ;
        RECT 66.200 14.800 70.600 15.100 ;
        RECT 90.200 14.800 90.600 15.200 ;
        RECT 91.000 15.100 91.400 15.200 ;
        RECT 134.200 15.100 134.600 15.200 ;
        RECT 149.400 15.100 149.800 15.200 ;
        RECT 91.000 14.800 149.800 15.100 ;
        RECT 6.200 14.100 6.600 14.200 ;
        RECT 19.000 14.100 19.400 14.200 ;
        RECT 6.200 13.800 19.400 14.100 ;
        RECT 24.600 14.100 25.000 14.200 ;
        RECT 26.200 14.100 26.600 14.200 ;
        RECT 24.600 13.800 26.600 14.100 ;
        RECT 30.200 14.100 30.600 14.200 ;
        RECT 31.800 14.100 32.200 14.200 ;
        RECT 30.200 13.800 32.200 14.100 ;
        RECT 38.200 14.100 38.600 14.200 ;
        RECT 40.600 14.100 41.000 14.200 ;
        RECT 38.200 13.800 41.000 14.100 ;
        RECT 46.200 14.100 46.600 14.200 ;
        RECT 51.000 14.100 51.400 14.200 ;
        RECT 46.200 13.800 51.400 14.100 ;
        RECT 72.600 14.100 73.000 14.200 ;
        RECT 76.600 14.100 77.000 14.200 ;
        RECT 72.600 13.800 77.000 14.100 ;
        RECT 90.200 14.100 90.500 14.800 ;
        RECT 99.000 14.100 99.400 14.200 ;
        RECT 105.400 14.100 105.800 14.200 ;
        RECT 90.200 13.800 105.800 14.100 ;
        RECT 106.200 14.100 106.600 14.200 ;
        RECT 110.200 14.100 110.600 14.200 ;
        RECT 106.200 13.800 110.600 14.100 ;
        RECT 111.000 14.100 111.400 14.200 ;
        RECT 128.600 14.100 129.000 14.200 ;
        RECT 136.600 14.100 137.000 14.200 ;
        RECT 111.000 13.800 137.000 14.100 ;
        RECT 111.000 13.200 111.300 13.800 ;
        RECT 4.600 13.100 5.000 13.200 ;
        RECT 11.800 13.100 12.200 13.200 ;
        RECT 23.800 13.100 24.200 13.200 ;
        RECT 27.800 13.100 28.200 13.200 ;
        RECT 49.400 13.100 49.800 13.200 ;
        RECT 4.600 12.800 49.800 13.100 ;
        RECT 86.200 13.100 86.600 13.200 ;
        RECT 91.800 13.100 92.200 13.200 ;
        RECT 86.200 12.800 92.200 13.100 ;
        RECT 94.200 13.100 94.600 13.200 ;
        RECT 99.800 13.100 100.200 13.200 ;
        RECT 104.600 13.100 105.000 13.200 ;
        RECT 109.400 13.100 109.800 13.200 ;
        RECT 94.200 12.800 109.800 13.100 ;
        RECT 111.000 12.800 111.400 13.200 ;
        RECT 111.800 12.800 112.200 13.200 ;
        RECT 112.600 13.100 113.000 13.200 ;
        RECT 124.600 13.100 125.000 13.200 ;
        RECT 128.600 13.100 129.000 13.200 ;
        RECT 134.200 13.100 134.600 13.200 ;
        RECT 112.600 12.800 129.000 13.100 ;
        RECT 131.000 12.800 134.600 13.100 ;
        RECT 135.800 13.100 136.200 13.200 ;
        RECT 142.200 13.100 142.600 13.200 ;
        RECT 135.800 12.800 142.600 13.100 ;
        RECT 9.400 12.100 9.800 12.200 ;
        RECT 12.600 12.100 13.000 12.200 ;
        RECT 9.400 11.800 13.000 12.100 ;
        RECT 19.000 12.100 19.400 12.200 ;
        RECT 23.800 12.100 24.200 12.200 ;
        RECT 35.000 12.100 35.400 12.200 ;
        RECT 19.000 11.800 35.400 12.100 ;
        RECT 45.400 12.100 45.800 12.200 ;
        RECT 46.200 12.100 46.600 12.200 ;
        RECT 45.400 11.800 46.600 12.100 ;
        RECT 69.400 12.100 69.800 12.200 ;
        RECT 107.800 12.100 108.200 12.200 ;
        RECT 69.400 11.800 108.200 12.100 ;
        RECT 108.600 12.100 109.000 12.200 ;
        RECT 111.800 12.100 112.100 12.800 ;
        RECT 131.000 12.200 131.300 12.800 ;
        RECT 108.600 11.800 112.100 12.100 ;
        RECT 120.600 12.100 121.000 12.200 ;
        RECT 123.800 12.100 124.200 12.200 ;
        RECT 120.600 11.800 124.200 12.100 ;
        RECT 131.000 11.800 131.400 12.200 ;
        RECT 137.400 12.100 137.800 12.200 ;
        RECT 139.800 12.100 140.200 12.200 ;
        RECT 137.400 11.800 140.200 12.100 ;
        RECT 17.400 11.100 17.800 11.200 ;
        RECT 35.800 11.100 36.200 11.200 ;
        RECT 39.000 11.100 39.400 11.200 ;
        RECT 17.400 10.800 39.400 11.100 ;
        RECT 53.400 11.100 53.800 11.200 ;
        RECT 64.600 11.100 65.000 11.200 ;
        RECT 53.400 10.800 65.000 11.100 ;
        RECT 83.000 11.100 83.400 11.200 ;
        RECT 85.400 11.100 85.800 11.200 ;
        RECT 89.400 11.100 89.800 11.200 ;
        RECT 83.000 10.800 89.800 11.100 ;
        RECT 110.200 11.100 110.600 11.200 ;
        RECT 117.400 11.100 117.800 11.200 ;
        RECT 110.200 10.800 117.800 11.100 ;
        RECT 141.400 11.100 141.800 11.200 ;
        RECT 143.000 11.100 143.400 11.200 ;
        RECT 141.400 10.800 143.400 11.100 ;
        RECT 10.200 10.100 10.600 10.200 ;
        RECT 23.000 10.100 23.400 10.200 ;
        RECT 28.600 10.100 29.000 10.200 ;
        RECT 30.200 10.100 30.600 10.200 ;
        RECT 10.200 9.800 30.600 10.100 ;
        RECT 35.000 10.100 35.400 10.200 ;
        RECT 35.800 10.100 36.200 10.200 ;
        RECT 35.000 9.800 36.200 10.100 ;
        RECT 36.600 10.100 37.000 10.200 ;
        RECT 58.200 10.100 58.600 10.200 ;
        RECT 36.600 9.800 58.600 10.100 ;
        RECT 66.200 10.100 66.600 10.200 ;
        RECT 107.800 10.100 108.200 10.200 ;
        RECT 111.000 10.100 111.400 10.200 ;
        RECT 115.000 10.100 115.400 10.200 ;
        RECT 66.200 9.800 97.700 10.100 ;
        RECT 107.800 9.800 115.400 10.100 ;
        RECT 5.400 9.100 5.800 9.200 ;
        RECT 11.800 9.100 12.200 9.200 ;
        RECT 18.200 9.100 18.600 9.200 ;
        RECT 33.400 9.100 33.800 9.200 ;
        RECT 63.800 9.100 64.200 9.200 ;
        RECT 5.400 8.800 64.200 9.100 ;
        RECT 71.000 9.100 71.400 9.200 ;
        RECT 71.800 9.100 72.200 9.200 ;
        RECT 71.000 8.800 72.200 9.100 ;
        RECT 78.200 8.800 78.600 9.200 ;
        RECT 81.400 9.100 81.800 9.200 ;
        RECT 82.200 9.100 82.600 9.200 ;
        RECT 86.200 9.100 86.600 9.200 ;
        RECT 81.400 8.800 86.600 9.100 ;
        RECT 87.800 9.100 88.200 9.200 ;
        RECT 96.600 9.100 97.000 9.200 ;
        RECT 87.800 8.800 97.000 9.100 ;
        RECT 97.400 9.100 97.700 9.800 ;
        RECT 107.000 9.100 107.400 9.200 ;
        RECT 114.200 9.100 114.600 9.200 ;
        RECT 116.600 9.100 117.000 9.200 ;
        RECT 97.400 8.800 117.000 9.100 ;
        RECT 129.400 9.100 129.800 9.200 ;
        RECT 134.200 9.100 134.600 9.200 ;
        RECT 138.200 9.100 138.600 9.200 ;
        RECT 129.400 8.800 138.600 9.100 ;
        RECT 3.000 8.100 3.400 8.200 ;
        RECT 6.200 8.100 6.600 8.200 ;
        RECT 3.000 7.800 6.600 8.100 ;
        RECT 27.800 7.800 28.200 8.200 ;
        RECT 37.400 7.800 37.800 8.200 ;
        RECT 70.200 8.100 70.600 8.200 ;
        RECT 75.800 8.100 76.200 8.200 ;
        RECT 70.200 7.800 76.200 8.100 ;
        RECT 78.200 8.100 78.500 8.800 ;
        RECT 89.400 8.100 89.800 8.200 ;
        RECT 78.200 7.800 89.800 8.100 ;
        RECT 91.000 8.100 91.400 8.200 ;
        RECT 100.600 8.100 101.000 8.200 ;
        RECT 112.600 8.100 113.000 8.200 ;
        RECT 91.000 7.800 113.000 8.100 ;
        RECT 122.200 7.800 122.600 8.200 ;
        RECT 127.800 8.100 128.200 8.200 ;
        RECT 143.800 8.100 144.200 8.200 ;
        RECT 146.200 8.100 146.600 8.200 ;
        RECT 127.800 7.800 146.600 8.100 ;
        RECT 27.800 7.100 28.100 7.800 ;
        RECT 37.400 7.100 37.700 7.800 ;
        RECT 122.200 7.200 122.500 7.800 ;
        RECT 27.800 6.800 37.700 7.100 ;
        RECT 41.400 7.100 41.800 7.200 ;
        RECT 45.400 7.100 45.800 7.200 ;
        RECT 49.400 7.100 49.800 7.200 ;
        RECT 41.400 6.800 49.800 7.100 ;
        RECT 54.200 7.100 54.600 7.200 ;
        RECT 55.800 7.100 56.200 7.200 ;
        RECT 54.200 6.800 56.200 7.100 ;
        RECT 74.200 7.100 74.600 7.200 ;
        RECT 79.800 7.100 80.200 7.200 ;
        RECT 84.600 7.100 85.000 7.200 ;
        RECT 74.200 6.800 85.000 7.100 ;
        RECT 86.200 7.100 86.600 7.200 ;
        RECT 90.200 7.100 90.600 7.200 ;
        RECT 86.200 6.800 90.600 7.100 ;
        RECT 91.800 7.100 92.200 7.200 ;
        RECT 94.200 7.100 94.600 7.200 ;
        RECT 111.000 7.100 111.400 7.200 ;
        RECT 115.000 7.100 115.400 7.200 ;
        RECT 91.800 6.800 94.600 7.100 ;
        RECT 95.000 6.800 115.400 7.100 ;
        RECT 118.200 7.100 118.600 7.200 ;
        RECT 119.800 7.100 120.200 7.200 ;
        RECT 118.200 6.800 120.200 7.100 ;
        RECT 122.200 6.800 122.600 7.200 ;
        RECT 123.800 7.100 124.200 7.200 ;
        RECT 128.600 7.100 129.000 7.200 ;
        RECT 123.800 6.800 129.000 7.100 ;
        RECT 131.800 7.100 132.200 7.200 ;
        RECT 136.600 7.100 137.000 7.200 ;
        RECT 131.800 6.800 137.000 7.100 ;
        RECT 145.400 7.100 145.800 7.200 ;
        RECT 148.600 7.100 149.000 7.200 ;
        RECT 145.400 6.800 149.000 7.100 ;
        RECT 95.000 6.200 95.300 6.800 ;
        RECT 15.800 6.100 16.200 6.200 ;
        RECT 37.400 6.100 37.800 6.200 ;
        RECT 39.800 6.100 40.200 6.200 ;
        RECT 15.800 5.800 40.200 6.100 ;
        RECT 48.600 6.100 49.000 6.200 ;
        RECT 52.600 6.100 53.000 6.200 ;
        RECT 48.600 5.800 53.000 6.100 ;
        RECT 71.000 6.100 71.400 6.200 ;
        RECT 73.400 6.100 73.800 6.200 ;
        RECT 71.000 5.800 73.800 6.100 ;
        RECT 74.200 6.100 74.600 6.200 ;
        RECT 79.000 6.100 79.400 6.200 ;
        RECT 82.200 6.100 82.600 6.200 ;
        RECT 92.600 6.100 93.000 6.200 ;
        RECT 74.200 5.800 93.000 6.100 ;
        RECT 95.000 5.800 95.400 6.200 ;
        RECT 102.200 6.100 102.600 6.200 ;
        RECT 103.800 6.100 104.200 6.200 ;
        RECT 102.200 5.800 104.200 6.100 ;
        RECT 107.800 6.100 108.200 6.200 ;
        RECT 111.000 6.100 111.400 6.200 ;
        RECT 107.800 5.800 111.400 6.100 ;
        RECT 120.600 6.100 121.000 6.200 ;
        RECT 121.400 6.100 121.800 6.200 ;
        RECT 120.600 5.800 121.800 6.100 ;
        RECT 129.400 6.100 129.800 6.200 ;
        RECT 131.800 6.100 132.200 6.200 ;
        RECT 129.400 5.800 132.200 6.100 ;
        RECT 137.400 6.100 137.800 6.200 ;
        RECT 142.200 6.100 142.600 6.200 ;
        RECT 146.200 6.100 146.600 6.200 ;
        RECT 137.400 5.800 146.600 6.100 ;
        RECT 26.200 5.100 26.600 5.200 ;
        RECT 31.000 5.100 31.400 5.200 ;
        RECT 26.200 4.800 31.400 5.100 ;
        RECT 79.000 5.100 79.400 5.200 ;
        RECT 86.200 5.100 86.600 5.200 ;
        RECT 87.800 5.100 88.200 5.200 ;
        RECT 79.000 4.800 80.100 5.100 ;
        RECT 86.200 4.800 88.200 5.100 ;
        RECT 131.000 5.100 131.400 5.200 ;
        RECT 131.800 5.100 132.200 5.200 ;
        RECT 131.000 4.800 132.200 5.100 ;
        RECT 133.400 5.100 133.800 5.200 ;
        RECT 139.800 5.100 140.200 5.200 ;
        RECT 133.400 4.800 140.200 5.100 ;
      LAYER via3 ;
        RECT 65.400 126.800 65.800 127.200 ;
        RECT 87.000 124.800 87.400 125.200 ;
        RECT 40.600 123.800 41.000 124.200 ;
        RECT 42.200 123.800 42.600 124.200 ;
        RECT 32.600 121.800 33.000 122.200 ;
        RECT 112.600 120.800 113.000 121.200 ;
        RECT 23.800 117.800 24.200 118.200 ;
        RECT 120.600 117.800 121.000 118.200 ;
        RECT 4.600 116.800 5.000 117.200 ;
        RECT 14.200 115.800 14.600 116.200 ;
        RECT 109.400 114.800 109.800 115.200 ;
        RECT 119.800 114.800 120.200 115.200 ;
        RECT 55.800 111.800 56.200 112.200 ;
        RECT 15.800 106.800 16.200 107.200 ;
        RECT 32.600 106.800 33.000 107.200 ;
        RECT 88.600 106.800 89.000 107.200 ;
        RECT 38.200 105.800 38.600 106.200 ;
        RECT 93.400 105.800 93.800 106.200 ;
        RECT 65.400 104.800 65.800 105.200 ;
        RECT 31.000 103.800 31.400 104.200 ;
        RECT 122.200 102.800 122.600 103.200 ;
        RECT 6.200 96.800 6.600 97.200 ;
        RECT 23.800 95.800 24.200 96.200 ;
        RECT 52.600 94.800 53.000 95.200 ;
        RECT 37.400 93.800 37.800 94.200 ;
        RECT 55.000 93.800 55.400 94.200 ;
        RECT 73.400 93.800 73.800 94.200 ;
        RECT 94.200 92.800 94.600 93.200 ;
        RECT 103.800 92.800 104.200 93.200 ;
        RECT 4.600 91.800 5.000 92.200 ;
        RECT 65.400 90.800 65.800 91.200 ;
        RECT 113.400 89.800 113.800 90.200 ;
        RECT 56.600 87.800 57.000 88.200 ;
        RECT 63.800 87.800 64.200 88.200 ;
        RECT 7.800 86.800 8.200 87.200 ;
        RECT 40.600 86.800 41.000 87.200 ;
        RECT 123.800 86.800 124.200 87.200 ;
        RECT 32.600 85.800 33.000 86.200 ;
        RECT 39.800 83.800 40.200 84.200 ;
        RECT 135.800 83.800 136.200 84.200 ;
        RECT 139.000 82.800 139.400 83.200 ;
        RECT 17.400 81.800 17.800 82.200 ;
        RECT 110.200 79.800 110.600 80.200 ;
        RECT 73.400 78.800 73.800 79.200 ;
        RECT 80.600 77.800 81.000 78.200 ;
        RECT 87.800 76.800 88.200 77.200 ;
        RECT 92.600 76.800 93.000 77.200 ;
        RECT 6.200 75.800 6.600 76.200 ;
        RECT 94.200 75.800 94.600 76.200 ;
        RECT 98.200 75.800 98.600 76.200 ;
        RECT 136.600 75.800 137.000 76.200 ;
        RECT 7.000 74.800 7.400 75.200 ;
        RECT 71.800 74.800 72.200 75.200 ;
        RECT 61.400 73.800 61.800 74.200 ;
        RECT 17.400 72.800 17.800 73.200 ;
        RECT 84.600 72.800 85.000 73.200 ;
        RECT 100.600 72.800 101.000 73.200 ;
        RECT 70.200 71.800 70.600 72.200 ;
        RECT 104.600 71.800 105.000 72.200 ;
        RECT 77.400 70.800 77.800 71.200 ;
        RECT 105.400 70.800 105.800 71.200 ;
        RECT 125.400 69.800 125.800 70.200 ;
        RECT 81.400 68.800 81.800 69.200 ;
        RECT 69.400 67.800 69.800 68.200 ;
        RECT 104.600 66.800 105.000 67.200 ;
        RECT 118.200 64.800 118.600 65.200 ;
        RECT 101.400 63.800 101.800 64.200 ;
        RECT 133.400 63.800 133.800 64.200 ;
        RECT 82.200 61.800 82.600 62.200 ;
        RECT 111.800 61.800 112.200 62.200 ;
        RECT 132.600 61.800 133.000 62.200 ;
        RECT 81.400 59.800 81.800 60.200 ;
        RECT 124.600 59.800 125.000 60.200 ;
        RECT 89.400 57.800 89.800 58.200 ;
        RECT 11.000 56.800 11.400 57.200 ;
        RECT 69.400 56.800 69.800 57.200 ;
        RECT 126.200 56.800 126.600 57.200 ;
        RECT 76.600 55.800 77.000 56.200 ;
        RECT 111.000 55.800 111.400 56.200 ;
        RECT 41.400 54.800 41.800 55.200 ;
        RECT 54.200 54.800 54.600 55.200 ;
        RECT 99.800 54.800 100.200 55.200 ;
        RECT 107.800 54.800 108.200 55.200 ;
        RECT 121.400 54.800 121.800 55.200 ;
        RECT 123.800 54.800 124.200 55.200 ;
        RECT 68.600 53.800 69.000 54.200 ;
        RECT 79.800 53.800 80.200 54.200 ;
        RECT 91.800 52.800 92.200 53.200 ;
        RECT 77.400 51.800 77.800 52.200 ;
        RECT 98.200 50.800 98.600 51.200 ;
        RECT 83.800 49.800 84.200 50.200 ;
        RECT 97.400 48.800 97.800 49.200 ;
        RECT 141.400 48.800 141.800 49.200 ;
        RECT 50.200 47.800 50.600 48.200 ;
        RECT 91.000 47.800 91.400 48.200 ;
        RECT 103.000 47.800 103.400 48.200 ;
        RECT 149.400 47.800 149.800 48.200 ;
        RECT 89.400 46.800 89.800 47.200 ;
        RECT 100.600 46.800 101.000 47.200 ;
        RECT 135.800 46.800 136.200 47.200 ;
        RECT 39.000 45.800 39.400 46.200 ;
        RECT 76.600 45.800 77.000 46.200 ;
        RECT 128.600 45.800 129.000 46.200 ;
        RECT 107.800 44.800 108.200 45.200 ;
        RECT 50.200 43.800 50.600 44.200 ;
        RECT 71.800 43.800 72.200 44.200 ;
        RECT 75.800 41.800 76.200 42.200 ;
        RECT 69.400 39.800 69.800 40.200 ;
        RECT 55.000 38.800 55.400 39.200 ;
        RECT 59.000 37.800 59.400 38.200 ;
        RECT 107.000 37.800 107.400 38.200 ;
        RECT 143.800 35.800 144.200 36.200 ;
        RECT 64.600 34.800 65.000 35.200 ;
        RECT 36.600 33.800 37.000 34.200 ;
        RECT 126.200 33.800 126.600 34.200 ;
        RECT 111.800 32.800 112.200 33.200 ;
        RECT 7.800 30.800 8.200 31.200 ;
        RECT 84.600 30.800 85.000 31.200 ;
        RECT 60.600 29.800 61.000 30.200 ;
        RECT 46.200 28.800 46.600 29.200 ;
        RECT 85.400 28.800 85.800 29.200 ;
        RECT 109.400 28.800 109.800 29.200 ;
        RECT 117.400 28.800 117.800 29.200 ;
        RECT 125.400 28.800 125.800 29.200 ;
        RECT 50.200 27.800 50.600 28.200 ;
        RECT 109.400 27.800 109.800 28.200 ;
        RECT 27.000 26.800 27.400 27.200 ;
        RECT 41.400 26.800 41.800 27.200 ;
        RECT 73.400 26.800 73.800 27.200 ;
        RECT 91.000 26.800 91.400 27.200 ;
        RECT 95.000 26.800 95.400 27.200 ;
        RECT 106.200 26.800 106.600 27.200 ;
        RECT 108.600 26.800 109.000 27.200 ;
        RECT 112.600 26.800 113.000 27.200 ;
        RECT 57.400 25.800 57.800 26.200 ;
        RECT 75.000 24.800 75.400 25.200 ;
        RECT 54.200 23.800 54.600 24.200 ;
        RECT 82.200 23.800 82.600 24.200 ;
        RECT 93.400 23.800 93.800 24.200 ;
        RECT 139.000 22.800 139.400 23.200 ;
        RECT 74.200 21.800 74.600 22.200 ;
        RECT 107.800 20.800 108.200 21.200 ;
        RECT 95.800 17.800 96.200 18.200 ;
        RECT 121.400 17.800 121.800 18.200 ;
        RECT 92.600 16.800 93.000 17.200 ;
        RECT 126.200 16.800 126.600 17.200 ;
        RECT 76.600 15.800 77.000 16.200 ;
        RECT 106.200 15.800 106.600 16.200 ;
        RECT 108.600 15.800 109.000 16.200 ;
        RECT 122.200 15.800 122.600 16.200 ;
        RECT 148.600 15.800 149.000 16.200 ;
        RECT 134.200 14.800 134.600 15.200 ;
        RECT 128.600 13.800 129.000 14.200 ;
        RECT 124.600 12.800 125.000 13.200 ;
        RECT 35.000 11.800 35.400 12.200 ;
        RECT 123.800 11.800 124.200 12.200 ;
        RECT 35.800 9.800 36.200 10.200 ;
        RECT 71.800 8.800 72.200 9.200 ;
        RECT 89.400 7.800 89.800 8.200 ;
        RECT 94.200 6.800 94.600 7.200 ;
        RECT 111.000 6.800 111.400 7.200 ;
        RECT 73.400 5.800 73.800 6.200 ;
        RECT 121.400 5.800 121.800 6.200 ;
        RECT 87.800 4.800 88.200 5.200 ;
        RECT 131.800 4.800 132.200 5.200 ;
      LAYER metal4 ;
        RECT 39.800 128.100 40.200 128.200 ;
        RECT 39.800 127.800 40.900 128.100 ;
        RECT 40.600 124.200 40.900 127.800 ;
        RECT 41.400 127.800 41.800 128.200 ;
        RECT 40.600 123.800 41.000 124.200 ;
        RECT 41.400 124.100 41.700 127.800 ;
        RECT 65.400 127.100 65.800 127.200 ;
        RECT 66.200 127.100 66.600 127.200 ;
        RECT 65.400 126.800 66.600 127.100 ;
        RECT 73.400 127.100 73.800 127.200 ;
        RECT 74.200 127.100 74.600 127.200 ;
        RECT 73.400 126.800 74.600 127.100 ;
        RECT 89.400 126.800 89.800 127.200 ;
        RECT 87.000 124.800 87.400 125.200 ;
        RECT 42.200 124.100 42.600 124.200 ;
        RECT 41.400 123.800 42.600 124.100 ;
        RECT 32.600 121.800 33.000 122.200 ;
        RECT 23.800 117.800 24.200 118.200 ;
        RECT 4.600 116.800 5.000 117.200 ;
        RECT 2.200 114.800 2.600 115.200 ;
        RECT 2.200 113.200 2.500 114.800 ;
        RECT 2.200 112.800 2.600 113.200 ;
        RECT 0.600 104.800 1.000 105.200 ;
        RECT 0.600 69.200 0.900 104.800 ;
        RECT 2.200 103.200 2.500 112.800 ;
        RECT 2.200 102.800 2.600 103.200 ;
        RECT 4.600 92.200 4.900 116.800 ;
        RECT 14.200 115.800 14.600 116.200 ;
        RECT 6.200 96.800 6.600 97.200 ;
        RECT 4.600 91.800 5.000 92.200 ;
        RECT 6.200 76.200 6.500 96.800 ;
        RECT 14.200 91.200 14.500 115.800 ;
        RECT 15.800 106.800 16.200 107.200 ;
        RECT 15.800 91.200 16.100 106.800 ;
        RECT 23.800 96.200 24.100 117.800 ;
        RECT 32.600 110.200 32.900 121.800 ;
        RECT 55.800 111.800 56.200 112.200 ;
        RECT 32.600 109.800 33.000 110.200 ;
        RECT 32.600 107.100 33.000 107.200 ;
        RECT 33.400 107.100 33.800 107.200 ;
        RECT 32.600 106.800 33.800 107.100 ;
        RECT 37.400 106.100 37.800 106.200 ;
        RECT 38.200 106.100 38.600 106.200 ;
        RECT 37.400 105.800 38.600 106.100 ;
        RECT 46.200 106.100 46.600 106.200 ;
        RECT 47.000 106.100 47.400 106.200 ;
        RECT 46.200 105.800 47.400 106.100 ;
        RECT 55.800 104.200 56.100 111.800 ;
        RECT 63.000 105.100 63.400 105.200 ;
        RECT 63.000 104.800 64.100 105.100 ;
        RECT 31.000 104.100 31.400 104.200 ;
        RECT 31.800 104.100 32.200 104.200 ;
        RECT 31.000 103.800 32.200 104.100 ;
        RECT 41.400 104.100 41.800 104.200 ;
        RECT 42.200 104.100 42.600 104.200 ;
        RECT 41.400 103.800 42.600 104.100 ;
        RECT 55.800 103.800 56.200 104.200 ;
        RECT 23.800 95.800 24.200 96.200 ;
        RECT 52.600 94.800 53.000 95.200 ;
        RECT 37.400 94.100 37.800 94.200 ;
        RECT 36.600 93.800 37.800 94.100 ;
        RECT 39.000 93.800 39.400 94.200 ;
        RECT 14.200 90.800 14.600 91.200 ;
        RECT 15.800 90.800 16.200 91.200 ;
        RECT 7.800 87.100 8.200 87.200 ;
        RECT 7.000 86.800 8.200 87.100 ;
        RECT 6.200 75.800 6.600 76.200 ;
        RECT 7.000 75.200 7.300 86.800 ;
        RECT 32.600 85.800 33.000 86.200 ;
        RECT 32.600 85.200 32.900 85.800 ;
        RECT 32.600 84.800 33.000 85.200 ;
        RECT 17.400 82.100 17.800 82.200 ;
        RECT 16.600 81.800 17.800 82.100 ;
        RECT 7.000 74.800 7.400 75.200 ;
        RECT 0.600 68.800 1.000 69.200 ;
        RECT 16.600 64.200 16.900 81.800 ;
        RECT 17.400 79.800 17.800 80.200 ;
        RECT 17.400 73.200 17.700 79.800 ;
        RECT 18.200 74.100 18.600 74.200 ;
        RECT 19.000 74.100 19.400 74.200 ;
        RECT 18.200 73.800 19.400 74.100 ;
        RECT 23.000 74.100 23.400 74.200 ;
        RECT 23.800 74.100 24.200 74.200 ;
        RECT 23.000 73.800 24.200 74.100 ;
        RECT 17.400 72.800 17.800 73.200 ;
        RECT 36.600 72.200 36.900 93.800 ;
        RECT 39.000 85.200 39.300 93.800 ;
        RECT 52.600 92.200 52.900 94.800 ;
        RECT 55.000 93.800 55.400 94.200 ;
        RECT 52.600 91.800 53.000 92.200 ;
        RECT 40.600 87.100 41.000 87.200 ;
        RECT 39.800 86.800 41.000 87.100 ;
        RECT 39.000 84.800 39.400 85.200 ;
        RECT 36.600 71.800 37.000 72.200 ;
        RECT 39.000 71.200 39.300 84.800 ;
        RECT 39.800 84.200 40.100 86.800 ;
        RECT 40.600 85.100 41.000 85.200 ;
        RECT 41.400 85.100 41.800 85.200 ;
        RECT 40.600 84.800 41.800 85.100 ;
        RECT 45.400 84.800 45.800 85.200 ;
        RECT 39.800 83.800 40.200 84.200 ;
        RECT 39.000 70.800 39.400 71.200 ;
        RECT 39.800 69.200 40.100 83.800 ;
        RECT 45.400 73.200 45.700 84.800 ;
        RECT 52.600 74.200 52.900 91.800 ;
        RECT 52.600 73.800 53.000 74.200 ;
        RECT 45.400 72.800 45.800 73.200 ;
        RECT 55.000 71.200 55.300 93.800 ;
        RECT 63.800 88.200 64.100 104.800 ;
        RECT 65.400 104.800 65.800 105.200 ;
        RECT 65.400 91.200 65.700 104.800 ;
        RECT 87.000 99.200 87.300 124.800 ;
        RECT 89.400 111.200 89.700 126.800 ;
        RECT 147.800 124.800 148.200 125.200 ;
        RECT 112.600 120.800 113.000 121.200 ;
        RECT 112.600 115.200 112.900 120.800 ;
        RECT 120.600 117.800 121.000 118.200 ;
        RECT 109.400 114.800 109.800 115.200 ;
        RECT 112.600 114.800 113.000 115.200 ;
        RECT 119.800 114.800 120.200 115.200 ;
        RECT 89.400 110.800 89.800 111.200 ;
        RECT 87.800 107.100 88.200 107.200 ;
        RECT 88.600 107.100 89.000 107.200 ;
        RECT 87.800 106.800 89.000 107.100 ;
        RECT 93.400 105.800 93.800 106.200 ;
        RECT 87.000 98.800 87.400 99.200 ;
        RECT 73.400 93.800 73.800 94.200 ;
        RECT 77.400 93.800 77.800 94.200 ;
        RECT 65.400 90.800 65.800 91.200 ;
        RECT 56.600 87.800 57.000 88.200 ;
        RECT 63.800 87.800 64.200 88.200 ;
        RECT 56.600 85.200 56.900 87.800 ;
        RECT 56.600 84.800 57.000 85.200 ;
        RECT 73.400 79.200 73.700 93.800 ;
        RECT 77.400 81.200 77.700 93.800 ;
        RECT 81.400 81.800 81.800 82.200 ;
        RECT 77.400 80.800 77.800 81.200 ;
        RECT 73.400 78.800 73.800 79.200 ;
        RECT 80.600 77.800 81.000 78.200 ;
        RECT 71.800 74.800 72.200 75.200 ;
        RECT 61.400 74.100 61.800 74.200 ;
        RECT 60.600 73.800 61.800 74.100 ;
        RECT 59.000 72.800 59.400 73.200 ;
        RECT 55.000 70.800 55.400 71.200 ;
        RECT 39.800 68.800 40.200 69.200 ;
        RECT 27.000 65.800 27.400 66.200 ;
        RECT 16.600 63.800 17.000 64.200 ;
        RECT 11.000 57.100 11.400 57.200 ;
        RECT 10.200 56.800 11.400 57.100 ;
        RECT 8.600 45.800 9.000 46.200 ;
        RECT 8.600 36.200 8.900 45.800 ;
        RECT 10.200 44.200 10.500 56.800 ;
        RECT 10.200 43.800 10.600 44.200 ;
        RECT 7.800 35.800 8.200 36.200 ;
        RECT 8.600 35.800 9.000 36.200 ;
        RECT 2.200 35.100 2.600 35.200 ;
        RECT 3.000 35.100 3.400 35.200 ;
        RECT 2.200 34.800 3.400 35.100 ;
        RECT 7.800 31.200 8.100 35.800 ;
        RECT 9.400 35.100 9.800 35.200 ;
        RECT 10.200 35.100 10.600 35.200 ;
        RECT 9.400 34.800 10.600 35.100 ;
        RECT 7.800 30.800 8.200 31.200 ;
        RECT 27.000 27.200 27.300 65.800 ;
        RECT 55.000 60.800 55.400 61.200 ;
        RECT 54.200 57.800 54.600 58.200 ;
        RECT 54.200 55.200 54.500 57.800 ;
        RECT 41.400 54.800 41.800 55.200 ;
        RECT 54.200 54.800 54.600 55.200 ;
        RECT 39.000 46.100 39.400 46.200 ;
        RECT 39.800 46.100 40.200 46.200 ;
        RECT 39.000 45.800 40.200 46.100 ;
        RECT 41.400 42.200 41.700 54.800 ;
        RECT 50.200 48.100 50.600 48.200 ;
        RECT 51.000 48.100 51.400 48.200 ;
        RECT 50.200 47.800 51.400 48.100 ;
        RECT 44.600 46.800 45.000 47.200 ;
        RECT 44.600 46.200 44.900 46.800 ;
        RECT 44.600 45.800 45.000 46.200 ;
        RECT 45.400 45.800 45.800 46.200 ;
        RECT 41.400 41.800 41.800 42.200 ;
        RECT 36.600 33.800 37.000 34.200 ;
        RECT 27.000 26.800 27.400 27.200 ;
        RECT 35.000 21.800 35.400 22.200 ;
        RECT 35.000 12.200 35.300 21.800 ;
        RECT 35.000 11.800 35.400 12.200 ;
        RECT 35.000 10.100 35.300 11.800 ;
        RECT 36.600 10.200 36.900 33.800 ;
        RECT 41.400 27.200 41.700 41.800 ;
        RECT 41.400 26.800 41.800 27.200 ;
        RECT 45.400 16.200 45.700 45.800 ;
        RECT 50.200 44.200 50.500 47.800 ;
        RECT 50.200 43.800 50.600 44.200 ;
        RECT 50.200 40.800 50.600 41.200 ;
        RECT 46.200 28.800 46.600 29.200 ;
        RECT 45.400 15.800 45.800 16.200 ;
        RECT 45.400 12.100 45.800 12.200 ;
        RECT 46.200 12.100 46.500 28.800 ;
        RECT 50.200 28.200 50.500 40.800 ;
        RECT 50.200 27.800 50.600 28.200 ;
        RECT 54.200 24.200 54.500 54.800 ;
        RECT 55.000 39.200 55.300 60.800 ;
        RECT 55.000 38.800 55.400 39.200 ;
        RECT 59.000 38.200 59.300 72.800 ;
        RECT 60.600 64.200 60.900 73.800 ;
        RECT 70.200 72.100 70.600 72.200 ;
        RECT 69.400 71.800 70.600 72.100 ;
        RECT 68.600 68.800 69.000 69.200 ;
        RECT 60.600 63.800 61.000 64.200 ;
        RECT 68.600 54.200 68.900 68.800 ;
        RECT 69.400 68.200 69.700 71.800 ;
        RECT 69.400 67.800 69.800 68.200 ;
        RECT 69.400 57.200 69.700 67.800 ;
        RECT 69.400 56.800 69.800 57.200 ;
        RECT 60.600 53.800 61.000 54.200 ;
        RECT 68.600 53.800 69.000 54.200 ;
        RECT 60.600 38.200 60.900 53.800 ;
        RECT 69.400 51.200 69.700 56.800 ;
        RECT 71.800 55.200 72.100 74.800 ;
        RECT 77.400 70.800 77.800 71.200 ;
        RECT 76.600 55.800 77.000 56.200 ;
        RECT 71.800 54.800 72.200 55.200 ;
        RECT 69.400 50.800 69.800 51.200 ;
        RECT 70.200 48.100 70.600 48.200 ;
        RECT 71.000 48.100 71.400 48.200 ;
        RECT 70.200 47.800 71.400 48.100 ;
        RECT 69.400 46.800 69.800 47.200 ;
        RECT 64.600 42.800 65.000 43.200 ;
        RECT 59.000 37.800 59.400 38.200 ;
        RECT 60.600 37.800 61.000 38.200 ;
        RECT 60.600 30.200 60.900 37.800 ;
        RECT 64.600 35.200 64.900 42.800 ;
        RECT 69.400 40.200 69.700 46.800 ;
        RECT 76.600 46.200 76.900 55.800 ;
        RECT 77.400 52.200 77.700 70.800 ;
        RECT 79.800 53.800 80.200 54.200 ;
        RECT 79.800 53.200 80.100 53.800 ;
        RECT 79.800 52.800 80.200 53.200 ;
        RECT 77.400 51.800 77.800 52.200 ;
        RECT 76.600 45.800 77.000 46.200 ;
        RECT 71.800 43.800 72.200 44.200 ;
        RECT 69.400 39.800 69.800 40.200 ;
        RECT 64.600 34.800 65.000 35.200 ;
        RECT 70.200 35.100 70.600 35.200 ;
        RECT 71.000 35.100 71.400 35.200 ;
        RECT 70.200 34.800 71.400 35.100 ;
        RECT 60.600 29.800 61.000 30.200 ;
        RECT 57.400 26.100 57.800 26.200 ;
        RECT 58.200 26.100 58.600 26.200 ;
        RECT 57.400 25.800 58.600 26.100 ;
        RECT 54.200 23.800 54.600 24.200 ;
        RECT 45.400 11.800 46.500 12.100 ;
        RECT 35.800 10.100 36.200 10.200 ;
        RECT 35.000 9.800 36.200 10.100 ;
        RECT 36.600 9.800 37.000 10.200 ;
        RECT 71.800 9.200 72.100 43.800 ;
        RECT 75.800 41.800 76.200 42.200 ;
        RECT 73.400 34.800 73.800 35.200 ;
        RECT 73.400 27.200 73.700 34.800 ;
        RECT 74.200 32.800 74.600 33.200 ;
        RECT 73.400 26.800 73.800 27.200 ;
        RECT 74.200 22.200 74.500 32.800 ;
        RECT 75.000 31.800 75.400 32.200 ;
        RECT 75.000 25.200 75.300 31.800 ;
        RECT 75.800 26.200 76.100 41.800 ;
        RECT 75.800 25.800 76.200 26.200 ;
        RECT 76.600 26.100 77.000 26.200 ;
        RECT 77.400 26.100 77.700 51.800 ;
        RECT 79.000 47.100 79.400 47.200 ;
        RECT 79.800 47.100 80.200 47.200 ;
        RECT 79.000 46.800 80.200 47.100 ;
        RECT 80.600 46.200 80.900 77.800 ;
        RECT 81.400 69.200 81.700 81.800 ;
        RECT 87.800 80.800 88.200 81.200 ;
        RECT 87.800 77.200 88.100 80.800 ;
        RECT 87.800 76.800 88.200 77.200 ;
        RECT 92.600 77.100 93.000 77.200 ;
        RECT 91.800 76.800 93.000 77.100 ;
        RECT 84.600 73.100 85.000 73.200 ;
        RECT 83.800 72.800 85.000 73.100 ;
        RECT 81.400 68.800 81.800 69.200 ;
        RECT 81.400 67.200 81.700 68.800 ;
        RECT 81.400 66.800 81.800 67.200 ;
        RECT 82.200 61.800 82.600 62.200 ;
        RECT 81.400 59.800 81.800 60.200 ;
        RECT 79.000 46.100 79.400 46.200 ;
        RECT 79.800 46.100 80.200 46.200 ;
        RECT 79.000 45.800 80.200 46.100 ;
        RECT 80.600 45.800 81.000 46.200 ;
        RECT 81.400 34.200 81.700 59.800 ;
        RECT 82.200 52.200 82.500 61.800 ;
        RECT 82.200 51.800 82.600 52.200 ;
        RECT 81.400 33.800 81.800 34.200 ;
        RECT 76.600 25.800 77.700 26.100 ;
        RECT 75.000 24.800 75.400 25.200 ;
        RECT 74.200 21.800 74.600 22.200 ;
        RECT 76.600 16.200 76.900 25.800 ;
        RECT 82.200 24.200 82.500 51.800 ;
        RECT 83.800 50.200 84.100 72.800 ;
        RECT 89.400 57.800 89.800 58.200 ;
        RECT 83.800 49.800 84.200 50.200 ;
        RECT 89.400 47.200 89.700 57.800 ;
        RECT 91.800 53.200 92.100 76.800 ;
        RECT 91.800 52.800 92.200 53.200 ;
        RECT 91.000 48.100 91.400 48.200 ;
        RECT 91.800 48.100 92.200 48.200 ;
        RECT 91.000 47.800 92.200 48.100 ;
        RECT 89.400 46.800 89.800 47.200 ;
        RECT 83.800 35.100 84.200 35.200 ;
        RECT 85.400 35.100 85.800 35.200 ;
        RECT 86.200 35.100 86.600 35.200 ;
        RECT 83.800 34.800 84.900 35.100 ;
        RECT 85.400 34.800 86.600 35.100 ;
        RECT 84.600 31.200 84.900 34.800 ;
        RECT 84.600 30.800 85.000 31.200 ;
        RECT 85.400 28.800 85.800 29.200 ;
        RECT 85.400 28.200 85.700 28.800 ;
        RECT 85.400 27.800 85.800 28.200 ;
        RECT 91.000 27.100 91.400 27.200 ;
        RECT 91.800 27.100 92.200 27.200 ;
        RECT 91.000 26.800 92.200 27.100 ;
        RECT 93.400 24.200 93.700 105.800 ;
        RECT 99.000 100.800 99.400 101.200 ;
        RECT 94.200 92.800 94.600 93.200 ;
        RECT 94.200 76.200 94.500 92.800 ;
        RECT 99.000 76.200 99.300 100.800 ;
        RECT 103.000 93.800 103.400 94.200 ;
        RECT 94.200 75.800 94.600 76.200 ;
        RECT 98.200 75.800 98.600 76.200 ;
        RECT 99.000 75.800 99.400 76.200 ;
        RECT 98.200 59.200 98.500 75.800 ;
        RECT 100.600 73.800 101.000 74.200 ;
        RECT 100.600 73.200 100.900 73.800 ;
        RECT 100.600 72.800 101.000 73.200 ;
        RECT 101.400 64.100 101.800 64.200 ;
        RECT 102.200 64.100 102.600 64.200 ;
        RECT 101.400 63.800 102.600 64.100 ;
        RECT 98.200 58.800 98.600 59.200 ;
        RECT 97.400 55.800 97.800 56.200 ;
        RECT 97.400 49.200 97.700 55.800 ;
        RECT 99.800 55.100 100.200 55.200 ;
        RECT 100.600 55.100 101.000 55.200 ;
        RECT 99.800 54.800 101.000 55.100 ;
        RECT 101.400 53.100 101.800 53.200 ;
        RECT 102.200 53.100 102.600 53.200 ;
        RECT 101.400 52.800 102.600 53.100 ;
        RECT 98.200 50.800 98.600 51.200 ;
        RECT 97.400 48.800 97.800 49.200 ;
        RECT 98.200 47.200 98.500 50.800 ;
        RECT 103.000 48.200 103.300 93.800 ;
        RECT 103.800 92.800 104.200 93.200 ;
        RECT 103.800 86.200 104.100 92.800 ;
        RECT 103.800 85.800 104.200 86.200 ;
        RECT 104.600 74.800 105.000 75.200 ;
        RECT 104.600 72.200 104.900 74.800 ;
        RECT 104.600 71.800 105.000 72.200 ;
        RECT 105.400 70.800 105.800 71.200 ;
        RECT 103.800 67.100 104.200 67.200 ;
        RECT 104.600 67.100 105.000 67.200 ;
        RECT 103.800 66.800 105.000 67.100 ;
        RECT 104.600 57.200 104.900 66.800 ;
        RECT 104.600 56.800 105.000 57.200 ;
        RECT 105.400 51.200 105.700 70.800 ;
        RECT 107.000 64.100 107.400 64.200 ;
        RECT 107.800 64.100 108.200 64.200 ;
        RECT 107.000 63.800 108.200 64.100 ;
        RECT 106.200 55.800 106.600 56.200 ;
        RECT 105.400 50.800 105.800 51.200 ;
        RECT 103.000 47.800 103.400 48.200 ;
        RECT 105.400 47.800 105.800 48.200 ;
        RECT 105.400 47.200 105.700 47.800 ;
        RECT 98.200 46.800 98.600 47.200 ;
        RECT 100.600 46.800 101.000 47.200 ;
        RECT 105.400 46.800 105.800 47.200 ;
        RECT 100.600 46.200 100.900 46.800 ;
        RECT 100.600 45.800 101.000 46.200 ;
        RECT 95.800 29.800 96.200 30.200 ;
        RECT 94.200 27.100 94.600 27.200 ;
        RECT 95.000 27.100 95.400 27.200 ;
        RECT 94.200 26.800 95.400 27.100 ;
        RECT 82.200 23.800 82.600 24.200 ;
        RECT 93.400 23.800 93.800 24.200 ;
        RECT 95.800 18.200 96.100 29.800 ;
        RECT 97.400 27.800 97.800 28.200 ;
        RECT 97.400 27.200 97.700 27.800 ;
        RECT 106.200 27.200 106.500 55.800 ;
        RECT 107.800 54.800 108.200 55.200 ;
        RECT 107.800 53.200 108.100 54.800 ;
        RECT 107.800 52.800 108.200 53.200 ;
        RECT 107.000 51.800 107.400 52.200 ;
        RECT 107.000 38.200 107.300 51.800 ;
        RECT 107.800 45.100 108.200 45.200 ;
        RECT 107.800 44.800 108.900 45.100 ;
        RECT 108.600 43.200 108.900 44.800 ;
        RECT 108.600 42.800 109.000 43.200 ;
        RECT 107.000 37.800 107.400 38.200 ;
        RECT 109.400 32.200 109.700 114.800 ;
        RECT 118.200 94.800 118.600 95.200 ;
        RECT 114.200 93.800 114.600 94.200 ;
        RECT 113.400 89.800 113.800 90.200 ;
        RECT 110.200 79.800 110.600 80.200 ;
        RECT 110.200 56.100 110.500 79.800 ;
        RECT 111.800 74.100 112.200 74.200 ;
        RECT 112.600 74.100 113.000 74.200 ;
        RECT 111.800 73.800 113.000 74.100 ;
        RECT 111.800 61.800 112.200 62.200 ;
        RECT 111.000 56.100 111.400 56.200 ;
        RECT 110.200 55.800 111.400 56.100 ;
        RECT 111.000 33.100 111.300 55.800 ;
        RECT 111.800 48.200 112.100 61.800 ;
        RECT 113.400 56.200 113.700 89.800 ;
        RECT 114.200 70.200 114.500 93.800 ;
        RECT 114.200 69.800 114.600 70.200 ;
        RECT 118.200 65.200 118.500 94.800 ;
        RECT 119.000 93.800 119.400 94.200 ;
        RECT 118.200 64.800 118.600 65.200 ;
        RECT 113.400 55.800 113.800 56.200 ;
        RECT 115.000 54.800 115.400 55.200 ;
        RECT 111.800 47.800 112.200 48.200 ;
        RECT 111.800 33.100 112.200 33.200 ;
        RECT 111.000 32.800 112.200 33.100 ;
        RECT 109.400 31.800 109.800 32.200 ;
        RECT 109.400 30.800 109.800 31.200 ;
        RECT 109.400 29.200 109.700 30.800 ;
        RECT 109.400 28.800 109.800 29.200 ;
        RECT 115.000 28.200 115.300 54.800 ;
        RECT 119.000 51.200 119.300 93.800 ;
        RECT 119.000 50.800 119.400 51.200 ;
        RECT 115.800 39.800 116.200 40.200 ;
        RECT 109.400 27.800 109.800 28.200 ;
        RECT 115.000 27.800 115.400 28.200 ;
        RECT 97.400 26.800 97.800 27.200 ;
        RECT 106.200 26.800 106.600 27.200 ;
        RECT 108.600 27.100 109.000 27.200 ;
        RECT 107.800 26.800 109.000 27.100 ;
        RECT 107.800 21.200 108.100 26.800 ;
        RECT 107.800 20.800 108.200 21.200 ;
        RECT 109.400 19.200 109.700 27.800 ;
        RECT 111.800 27.100 112.200 27.200 ;
        RECT 112.600 27.100 113.000 27.200 ;
        RECT 111.800 26.800 113.000 27.100 ;
        RECT 115.000 27.100 115.400 27.200 ;
        RECT 115.800 27.100 116.100 39.800 ;
        RECT 119.800 39.200 120.100 114.800 ;
        RECT 120.600 114.200 120.900 117.800 ;
        RECT 120.600 113.800 121.000 114.200 ;
        RECT 147.000 109.800 147.400 110.200 ;
        RECT 122.200 102.800 122.600 103.200 ;
        RECT 120.600 55.100 121.000 55.200 ;
        RECT 121.400 55.100 121.800 55.200 ;
        RECT 120.600 54.800 121.800 55.100 ;
        RECT 119.800 38.800 120.200 39.200 ;
        RECT 117.400 28.800 117.800 29.200 ;
        RECT 115.000 26.800 116.100 27.100 ;
        RECT 116.600 27.800 117.000 28.200 ;
        RECT 116.600 27.200 116.900 27.800 ;
        RECT 116.600 26.800 117.000 27.200 ;
        RECT 115.800 26.200 116.100 26.800 ;
        RECT 115.800 25.800 116.200 26.200 ;
        RECT 117.400 25.200 117.700 28.800 ;
        RECT 122.200 25.200 122.500 102.800 ;
        RECT 123.800 87.100 124.200 87.200 ;
        RECT 124.600 87.100 125.000 87.200 ;
        RECT 123.800 86.800 125.000 87.100 ;
        RECT 129.400 87.100 129.800 87.200 ;
        RECT 130.200 87.100 130.600 87.200 ;
        RECT 129.400 86.800 130.600 87.100 ;
        RECT 135.800 83.800 136.200 84.200 ;
        RECT 125.400 69.800 125.800 70.200 ;
        RECT 123.000 65.800 123.400 66.200 ;
        RECT 123.000 27.200 123.300 65.800 ;
        RECT 124.600 59.800 125.000 60.200 ;
        RECT 123.800 54.800 124.200 55.200 ;
        RECT 123.800 53.200 124.100 54.800 ;
        RECT 124.600 54.200 124.900 59.800 ;
        RECT 124.600 53.800 125.000 54.200 ;
        RECT 123.800 52.800 124.200 53.200 ;
        RECT 124.600 50.200 124.900 53.800 ;
        RECT 124.600 49.800 125.000 50.200 ;
        RECT 123.000 27.100 123.400 27.200 ;
        RECT 123.000 26.800 124.100 27.100 ;
        RECT 117.400 24.800 117.800 25.200 ;
        RECT 122.200 24.800 122.600 25.200 ;
        RECT 109.400 18.800 109.800 19.200 ;
        RECT 95.800 17.800 96.200 18.200 ;
        RECT 121.400 17.800 121.800 18.200 ;
        RECT 92.600 17.100 93.000 17.200 ;
        RECT 93.400 17.100 93.800 17.200 ;
        RECT 92.600 16.800 93.800 17.100 ;
        RECT 76.600 15.800 77.000 16.200 ;
        RECT 106.200 15.800 106.600 16.200 ;
        RECT 108.600 15.800 109.000 16.200 ;
        RECT 106.200 14.200 106.500 15.800 ;
        RECT 106.200 13.800 106.600 14.200 ;
        RECT 108.600 12.200 108.900 15.800 ;
        RECT 111.000 13.800 111.400 14.200 ;
        RECT 108.600 11.800 109.000 12.200 ;
        RECT 71.800 8.800 72.200 9.200 ;
        RECT 87.800 8.800 88.200 9.200 ;
        RECT 74.200 6.800 74.600 7.200 ;
        RECT 73.400 6.100 73.800 6.200 ;
        RECT 74.200 6.100 74.500 6.800 ;
        RECT 73.400 5.800 74.500 6.100 ;
        RECT 87.800 5.200 88.100 8.800 ;
        RECT 89.400 8.100 89.800 8.200 ;
        RECT 90.200 8.100 90.600 8.200 ;
        RECT 89.400 7.800 90.600 8.100 ;
        RECT 111.000 7.200 111.300 13.800 ;
        RECT 94.200 6.800 94.600 7.200 ;
        RECT 111.000 6.800 111.400 7.200 ;
        RECT 94.200 5.200 94.500 6.800 ;
        RECT 121.400 6.200 121.700 17.800 ;
        RECT 122.200 16.800 122.600 17.200 ;
        RECT 122.200 16.200 122.500 16.800 ;
        RECT 122.200 15.800 122.600 16.200 ;
        RECT 122.200 7.200 122.500 15.800 ;
        RECT 123.800 12.200 124.100 26.800 ;
        RECT 124.600 13.200 124.900 49.800 ;
        RECT 125.400 41.200 125.700 69.800 ;
        RECT 133.400 64.100 133.800 64.200 ;
        RECT 132.600 63.800 133.800 64.100 ;
        RECT 132.600 62.200 132.900 63.800 ;
        RECT 132.600 61.800 133.000 62.200 ;
        RECT 126.200 56.800 126.600 57.200 ;
        RECT 126.200 52.200 126.500 56.800 ;
        RECT 126.200 51.800 126.600 52.200 ;
        RECT 126.200 47.800 126.600 48.200 ;
        RECT 128.600 47.800 129.000 48.200 ;
        RECT 125.400 40.800 125.800 41.200 ;
        RECT 126.200 34.200 126.500 47.800 ;
        RECT 128.600 47.200 128.900 47.800 ;
        RECT 128.600 46.800 129.000 47.200 ;
        RECT 128.600 46.200 128.900 46.800 ;
        RECT 128.600 45.800 129.000 46.200 ;
        RECT 132.600 40.200 132.900 61.800 ;
        RECT 133.400 55.800 133.800 56.200 ;
        RECT 133.400 55.200 133.700 55.800 ;
        RECT 133.400 54.800 133.800 55.200 ;
        RECT 135.800 47.200 136.100 83.800 ;
        RECT 139.000 82.800 139.400 83.200 ;
        RECT 139.000 76.200 139.300 82.800 ;
        RECT 136.600 75.800 137.000 76.200 ;
        RECT 139.000 75.800 139.400 76.200 ;
        RECT 134.200 46.800 134.600 47.200 ;
        RECT 135.800 46.800 136.200 47.200 ;
        RECT 132.600 39.800 133.000 40.200 ;
        RECT 126.200 33.800 126.600 34.200 ;
        RECT 126.200 29.200 126.500 33.800 ;
        RECT 128.600 32.800 129.000 33.200 ;
        RECT 125.400 28.800 125.800 29.200 ;
        RECT 126.200 28.800 126.600 29.200 ;
        RECT 125.400 27.200 125.700 28.800 ;
        RECT 125.400 26.800 125.800 27.200 ;
        RECT 126.200 20.800 126.600 21.200 ;
        RECT 126.200 17.200 126.500 20.800 ;
        RECT 126.200 16.800 126.600 17.200 ;
        RECT 127.000 17.100 127.400 17.200 ;
        RECT 127.800 17.100 128.200 17.200 ;
        RECT 127.000 16.800 128.200 17.100 ;
        RECT 128.600 14.200 128.900 32.800 ;
        RECT 133.400 19.800 133.800 20.200 ;
        RECT 133.400 19.200 133.700 19.800 ;
        RECT 133.400 18.800 133.800 19.200 ;
        RECT 134.200 15.200 134.500 46.800 ;
        RECT 136.600 46.200 136.900 75.800 ;
        RECT 136.600 45.800 137.000 46.200 ;
        RECT 139.000 23.200 139.300 75.800 ;
        RECT 141.400 71.800 141.800 72.200 ;
        RECT 141.400 49.200 141.700 71.800 ;
        RECT 143.800 63.800 144.200 64.200 ;
        RECT 141.400 48.800 141.800 49.200 ;
        RECT 143.800 36.200 144.100 63.800 ;
        RECT 147.000 53.200 147.300 109.800 ;
        RECT 147.000 52.800 147.400 53.200 ;
        RECT 147.800 49.200 148.100 124.800 ;
        RECT 148.600 93.800 149.000 94.200 ;
        RECT 148.600 55.200 148.900 93.800 ;
        RECT 148.600 54.800 149.000 55.200 ;
        RECT 147.800 48.800 148.200 49.200 ;
        RECT 143.800 35.800 144.200 36.200 ;
        RECT 139.000 22.800 139.400 23.200 ;
        RECT 148.600 16.200 148.900 54.800 ;
        RECT 149.400 50.800 149.800 51.200 ;
        RECT 149.400 48.200 149.700 50.800 ;
        RECT 149.400 47.800 149.800 48.200 ;
        RECT 148.600 15.800 149.000 16.200 ;
        RECT 134.200 14.800 134.600 15.200 ;
        RECT 128.600 13.800 129.000 14.200 ;
        RECT 124.600 12.800 125.000 13.200 ;
        RECT 123.800 11.800 124.200 12.200 ;
        RECT 127.000 8.100 127.400 8.200 ;
        RECT 127.800 8.100 128.200 8.200 ;
        RECT 127.000 7.800 128.200 8.100 ;
        RECT 122.200 6.800 122.600 7.200 ;
        RECT 131.800 6.800 132.200 7.200 ;
        RECT 121.400 5.800 121.800 6.200 ;
        RECT 131.800 5.200 132.100 6.800 ;
        RECT 87.800 4.800 88.200 5.200 ;
        RECT 94.200 4.800 94.600 5.200 ;
        RECT 131.000 5.100 131.400 5.200 ;
        RECT 131.800 5.100 132.200 5.200 ;
        RECT 131.000 4.800 132.200 5.100 ;
      LAYER via4 ;
        RECT 66.200 126.800 66.600 127.200 ;
        RECT 74.200 126.800 74.600 127.200 ;
        RECT 33.400 106.800 33.800 107.200 ;
        RECT 31.800 103.800 32.200 104.200 ;
        RECT 19.000 73.800 19.400 74.200 ;
        RECT 3.000 34.800 3.400 35.200 ;
        RECT 39.800 45.800 40.200 46.200 ;
        RECT 51.000 47.800 51.400 48.200 ;
        RECT 71.000 34.800 71.400 35.200 ;
        RECT 58.200 25.800 58.600 26.200 ;
        RECT 79.800 45.800 80.200 46.200 ;
        RECT 91.800 47.800 92.200 48.200 ;
        RECT 91.800 26.800 92.200 27.200 ;
        RECT 102.200 63.800 102.600 64.200 ;
        RECT 100.600 54.800 101.000 55.200 ;
        RECT 124.600 86.800 125.000 87.200 ;
        RECT 93.400 16.800 93.800 17.200 ;
        RECT 90.200 7.800 90.600 8.200 ;
      LAYER metal5 ;
        RECT 66.200 127.100 66.600 127.200 ;
        RECT 74.200 127.100 74.600 127.200 ;
        RECT 66.200 126.800 74.600 127.100 ;
        RECT 33.400 107.100 33.800 107.200 ;
        RECT 87.800 107.100 88.200 107.200 ;
        RECT 33.400 106.800 88.200 107.100 ;
        RECT 37.400 106.100 37.800 106.200 ;
        RECT 46.200 106.100 46.600 106.200 ;
        RECT 37.400 105.800 46.600 106.100 ;
        RECT 31.800 104.100 32.200 104.200 ;
        RECT 41.400 104.100 41.800 104.200 ;
        RECT 31.800 103.800 41.800 104.100 ;
        RECT 124.600 87.100 125.000 87.200 ;
        RECT 129.400 87.100 129.800 87.200 ;
        RECT 124.600 86.800 129.800 87.100 ;
        RECT 32.600 85.100 33.000 85.200 ;
        RECT 40.600 85.100 41.000 85.200 ;
        RECT 32.600 84.800 41.000 85.100 ;
        RECT 19.000 74.100 19.400 74.200 ;
        RECT 23.000 74.100 23.400 74.200 ;
        RECT 19.000 73.800 23.400 74.100 ;
        RECT 100.600 74.100 101.000 74.200 ;
        RECT 111.800 74.100 112.200 74.200 ;
        RECT 100.600 73.800 112.200 74.100 ;
        RECT 81.400 67.100 81.800 67.200 ;
        RECT 103.800 67.100 104.200 67.200 ;
        RECT 81.400 66.800 104.200 67.100 ;
        RECT 102.200 64.100 102.600 64.200 ;
        RECT 107.000 64.100 107.400 64.200 ;
        RECT 102.200 63.800 107.400 64.100 ;
        RECT 97.400 56.100 97.800 56.200 ;
        RECT 97.400 55.800 133.700 56.100 ;
        RECT 133.400 55.200 133.700 55.800 ;
        RECT 100.600 55.100 101.000 55.200 ;
        RECT 120.600 55.100 121.000 55.200 ;
        RECT 100.600 54.800 121.000 55.100 ;
        RECT 133.400 54.800 133.800 55.200 ;
        RECT 79.800 53.100 80.200 53.200 ;
        RECT 101.400 53.100 101.800 53.200 ;
        RECT 123.800 53.100 124.200 53.200 ;
        RECT 79.800 52.800 124.200 53.100 ;
        RECT 51.000 48.100 51.400 48.200 ;
        RECT 70.200 48.100 70.600 48.200 ;
        RECT 51.000 47.800 70.600 48.100 ;
        RECT 91.800 48.100 92.200 48.200 ;
        RECT 105.400 48.100 105.800 48.200 ;
        RECT 91.800 47.800 105.800 48.100 ;
        RECT 69.400 47.100 69.800 47.200 ;
        RECT 79.000 47.100 79.400 47.200 ;
        RECT 69.400 46.800 79.400 47.100 ;
        RECT 98.200 47.100 98.600 47.200 ;
        RECT 128.600 47.100 129.000 47.200 ;
        RECT 98.200 46.800 129.000 47.100 ;
        RECT 39.800 46.100 40.200 46.200 ;
        RECT 44.600 46.100 45.000 46.200 ;
        RECT 39.800 45.800 45.000 46.100 ;
        RECT 79.800 46.100 80.200 46.200 ;
        RECT 100.600 46.100 101.000 46.200 ;
        RECT 79.800 45.800 101.000 46.100 ;
        RECT 64.600 43.100 65.000 43.200 ;
        RECT 108.600 43.100 109.000 43.200 ;
        RECT 64.600 42.800 109.000 43.100 ;
        RECT 3.000 35.100 3.400 35.200 ;
        RECT 9.400 35.100 9.800 35.200 ;
        RECT 3.000 34.800 9.800 35.100 ;
        RECT 71.000 35.100 71.400 35.200 ;
        RECT 85.400 35.100 85.800 35.200 ;
        RECT 71.000 34.800 85.800 35.100 ;
        RECT 85.400 28.100 85.800 28.200 ;
        RECT 97.400 28.100 97.800 28.200 ;
        RECT 115.000 28.100 115.400 28.200 ;
        RECT 85.400 27.800 115.400 28.100 ;
        RECT 116.600 27.800 117.000 28.200 ;
        RECT 91.800 27.100 92.200 27.200 ;
        RECT 94.200 27.100 94.600 27.200 ;
        RECT 91.800 26.800 94.600 27.100 ;
        RECT 111.800 27.100 112.200 27.200 ;
        RECT 116.600 27.100 116.900 27.800 ;
        RECT 111.800 26.800 116.900 27.100 ;
        RECT 58.200 26.100 58.600 26.200 ;
        RECT 115.800 26.100 116.200 26.200 ;
        RECT 58.200 25.800 116.200 26.100 ;
        RECT 109.400 19.100 109.800 19.200 ;
        RECT 133.400 19.100 133.800 19.200 ;
        RECT 109.400 18.800 133.800 19.100 ;
        RECT 93.400 17.100 93.800 17.200 ;
        RECT 122.200 17.100 122.600 17.200 ;
        RECT 127.000 17.100 127.400 17.200 ;
        RECT 93.400 16.800 127.400 17.100 ;
        RECT 90.200 8.100 90.600 8.200 ;
        RECT 127.000 8.100 127.400 8.200 ;
        RECT 90.200 7.800 127.400 8.100 ;
        RECT 94.200 5.100 94.600 5.200 ;
        RECT 131.000 5.100 131.400 5.200 ;
        RECT 94.200 4.800 131.400 5.100 ;
  END
END alu
END LIBRARY

