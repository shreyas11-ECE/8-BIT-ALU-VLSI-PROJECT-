* NGSPICE file created from alu.ext - technology: scmos

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

.subckt alu vdd gnd a[0] a[1] a[2] a[3] a[4] a[5] a[6] a[7] b[0] b[1] b[2] b[3] b[4]
+ b[5] b[6] b[7] clk rst en opcode[0] opcode[1] opcode[2] out[0] out[1] out[2] out[3]
+ out[4] out[5] out[6] out[7] zero
XAND2X2_5 AND2X2_5/A a[7] gnd AND2X2_5/Y vdd AND2X2
XNAND2X1_10 NAND3X1_82/A NAND3X1_77/Y gnd NAND2X1_10/Y vdd NAND2X1
XNAND2X1_43 INVX2_16/Y INVX1_30/A gnd AOI21X1_38/A vdd NAND2X1
XNAND2X1_32 INVX8_2/Y MUX2X1_1/A gnd OAI21X1_9/B vdd NAND2X1
XNAND2X1_65 BUFX4_13/Y a[5] gnd NOR2X1_71/B vdd NAND2X1
XNAND2X1_21 NAND2X1_21/A NAND2X1_21/B gnd AOI21X1_25/C vdd NAND2X1
XNAND2X1_54 a[2] b[3] gnd OAI22X1_3/A vdd NAND2X1
XOAI22X1_3 OAI22X1_3/A OAI22X1_3/B AND2X2_13/Y INVX1_42/A gnd OR2X2_1/A vdd OAI22X1
XINVX2_12 INVX2_12/A gnd INVX2_12/Y vdd INVX2
XINVX2_23 OR2X2_9/B gnd INVX2_23/Y vdd INVX2
XFILL_11_1_0 gnd vdd FILL
XOAI21X1_19 OAI21X1_19/A OAI21X1_19/B AND2X2_4/Y gnd NAND3X1_19/C vdd OAI21X1
XFILL_12_3 gnd vdd FILL
XXNOR2X1_6 XNOR2X1_6/A INVX1_25/Y gnd NOR2X1_44/B vdd XNOR2X1
XFILL_0_0_0 gnd vdd FILL
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XOR2X2_11 OR2X2_11/A OR2X2_11/B gnd OR2X2_11/Y vdd OR2X2
XOR2X2_4 OR2X2_4/A INVX2_5/Y gnd OR2X2_4/Y vdd OR2X2
XFILL_8_1_0 gnd vdd FILL
XAND2X2_6 AND2X2_6/A AND2X2_6/B gnd AND2X2_6/Y vdd AND2X2
XAOI22X1_1 AOI22X1_1/A AOI22X1_1/B AOI22X1_1/C AOI22X1_1/D gnd AOI22X1_1/Y vdd AOI22X1
XNAND2X1_11 AOI22X1_1/B AOI22X1_1/A gnd AOI21X1_19/C vdd NAND2X1
XNAND2X1_55 NAND3X1_45/Y NAND2X1_55/B gnd NAND3X1_48/A vdd NAND2X1
XNAND2X1_22 BUFX4_3/Y a[2] gnd NOR2X1_47/B vdd NAND2X1
XNAND2X1_44 INVX8_2/Y AND2X2_5/Y gnd NOR2X1_15/A vdd NAND2X1
XNAND2X1_66 BUFX4_9/Y a[4] gnd INVX1_43/A vdd NAND2X1
XNAND2X1_33 NOR2X1_50/A INVX2_11/Y gnd OAI21X1_63/C vdd NAND2X1
XOAI22X1_4 NOR2X1_61/A NAND2X1_7/Y OAI22X1_4/C INVX1_43/A gnd INVX1_6/A vdd OAI22X1
XINVX2_13 en gnd INVX2_13/Y vdd INVX2
XFILL_11_1_1 gnd vdd FILL
XINVX2_24 b[6] gnd NOR2X1_7/B vdd INVX2
XFILL_10_1 gnd vdd FILL
XXNOR2X1_7 OR2X2_6/Y INVX2_16/Y gnd XNOR2X1_7/Y vdd XNOR2X1
XOR2X2_5 OR2X2_5/A OR2X2_5/B gnd OR2X2_5/Y vdd OR2X2
XFILL_0_0_1 gnd vdd FILL
XFILL_8_1_1 gnd vdd FILL
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XAND2X2_7 AND2X2_7/A AND2X2_7/B gnd AND2X2_7/Y vdd AND2X2
XNAND2X1_12 INVX2_2/Y NOR2X1_11/B gnd NAND2X1_12/Y vdd NAND2X1
XNAND2X1_34 NOR2X1_46/Y NOR2X1_45/Y gnd NAND2X1_34/Y vdd NAND2X1
XAOI22X1_2 INVX1_24/A AOI22X1_2/B AND2X2_8/Y INVX1_21/Y gnd AOI22X1_2/Y vdd AOI22X1
XNAND2X1_23 INVX8_2/A AND2X2_5/Y gnd NAND2X1_23/Y vdd NAND2X1
XNAND2X1_56 NOR2X1_5/A a[4] gnd OAI22X1_8/B vdd NAND2X1
XNAND2X1_67 BUFX4_1/Y a[6] gnd NOR2X1_71/A vdd NAND2X1
XNAND2X1_45 INVX8_2/Y INVX1_40/A gnd OAI21X1_73/C vdd NAND2X1
XAOI22X1_10 BUFX4_2/Y a[6] BUFX4_14/Y a[5] gnd OAI22X1_4/C vdd AOI22X1
XOAI22X1_5 OR2X2_4/Y OR2X2_2/B INVX4_5/Y OAI22X1_5/D gnd NOR2X1_16/B vdd OAI22X1
XINVX2_14 INVX2_14/A gnd INVX2_14/Y vdd INVX2
XINVX2_25 XOR2X1_5/Y gnd INVX2_25/Y vdd INVX2
XINVX8_1 rst gnd DFFSR_6/R vdd INVX8
XBUFX4_10 b[1] gnd NOR2X1_5/A vdd BUFX4
XOR2X2_6 OR2X2_6/A OR2X2_6/B gnd OR2X2_6/Y vdd OR2X2
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XAND2X2_8 AND2X2_8/A AND2X2_8/B gnd AND2X2_8/Y vdd AND2X2
XAOI22X1_3 INVX4_7/A INVX1_23/Y INVX2_11/Y AND2X2_6/Y gnd AOI22X1_3/Y vdd AOI22X1
XAOI22X1_11 NOR3X1_5/C NOR2X1_72/Y NOR2X1_11/B AOI22X1_11/D gnd AOI22X1_11/Y vdd AOI22X1
XNAND2X1_13 INVX2_2/A NOR2X1_11/B gnd AOI22X1_1/C vdd NAND2X1
XNAND2X1_35 a[0] b[3] gnd INVX2_14/A vdd NAND2X1
XNAND2X1_46 a[1] b[4] gnd OAI21X1_76/B vdd NAND2X1
XNAND2X1_68 NAND2X1_68/A NAND2X1_68/B gnd OAI21X1_18/B vdd NAND2X1
XNOR3X1_1 NOR3X1_1/A INVX1_7/A NOR3X1_1/C gnd NOR3X1_1/Y vdd NOR3X1
XNAND2X1_57 BUFX4_7/Y a[3] gnd INVX2_20/A vdd NAND2X1
XNAND2X1_24 BUFX4_7/Y NAND2X1_24/B gnd NAND2X1_24/Y vdd NAND2X1
XOAI22X1_6 NOR2X1_47/B OAI22X1_6/B AND2X2_9/Y INVX2_15/A gnd OAI22X1_6/Y vdd OAI22X1
XINVX2_15 INVX2_15/A gnd INVX2_15/Y vdd INVX2
XFILL_3_0_0 gnd vdd FILL
XINVX8_2 INVX8_2/A gnd INVX8_2/Y vdd INVX8
XBUFX4_11 b[1] gnd BUFX4_11/Y vdd BUFX4
XOR2X2_7 OR2X2_7/A OR2X2_7/B gnd OR2X2_7/Y vdd OR2X2
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XAND2X2_9 AND2X2_9/A AND2X2_9/B gnd AND2X2_9/Y vdd AND2X2
XAOI22X1_4 INVX2_11/Y INVX2_16/Y INVX4_5/A INVX1_29/Y gnd AOI22X1_4/Y vdd AOI22X1
XNAND2X1_36 INVX4_1/A a[1] gnd INVX2_15/A vdd NAND2X1
XNAND2X1_58 NAND2X1_58/A NAND2X1_58/B gnd NAND3X1_54/A vdd NAND2X1
XNAND2X1_47 a[1] b[3] gnd NOR2X1_60/B vdd NAND2X1
XNAND2X1_14 a[7] b[7] gnd INVX1_9/A vdd NAND2X1
XNOR3X1_2 INVX1_6/A NOR3X1_3/B NOR3X1_1/Y gnd NOR3X1_2/Y vdd NOR3X1
XNAND2X1_25 a[1] BUFX4_14/Y gnd AND2X2_6/B vdd NAND2X1
XOAI22X1_7 OR2X2_4/Y NOR2X1_3/A INVX4_5/Y NOR2X1_55/Y gnd NOR2X1_59/B vdd OAI22X1
XINVX2_16 INVX2_16/A gnd INVX2_16/Y vdd INVX2
XFILL_3_0_1 gnd vdd FILL
XBUFX4_12 b[1] gnd INVX8_2/A vdd BUFX4
XOR2X2_8 OR2X2_8/A OR2X2_8/B gnd OR2X2_8/Y vdd OR2X2
XAOI22X1_5 INVX1_12/Y INVX2_13/Y AOI22X1_5/C AOI22X1_5/D gnd DFFSR_4/D vdd AOI22X1
XNAND2X1_59 OR2X2_9/B OR2X2_9/A gnd NAND2X1_59/Y vdd NAND2X1
XNAND2X1_15 BUFX4_4/Y a[5] gnd NOR2X1_61/A vdd NAND2X1
XNAND2X1_48 BUFX4_5/Y a[4] gnd NOR2X1_52/A vdd NAND2X1
XNAND2X1_37 BUFX4_2/Y a[3] gnd AND2X2_9/A vdd NAND2X1
XNAND2X1_26 INVX2_10/Y INVX8_2/Y gnd AND2X2_6/A vdd NAND2X1
XNOR3X1_3 AND2X2_3/Y NOR3X1_3/B NOR3X1_1/Y gnd NOR3X1_3/Y vdd NOR3X1
XOAI22X1_8 AND2X2_9/A OAI22X1_8/B OAI22X1_8/C INVX2_12/A gnd INVX2_21/A vdd OAI22X1
XINVX2_17 b[4] gnd INVX2_17/Y vdd INVX2
XMUX2X1_1 MUX2X1_1/A MUX2X1_1/B BUFX4_11/Y gnd INVX1_14/A vdd MUX2X1
XBUFX4_13 b[1] gnd BUFX4_13/Y vdd BUFX4
XOR2X2_9 OR2X2_9/A OR2X2_9/B gnd OR2X2_9/Y vdd OR2X2
XFILL_7_1 gnd vdd FILL
XFILL_1_1_0 gnd vdd FILL
XNAND3X1_1 a[4] INVX2_17/Y INVX2_23/Y gnd OAI21X1_1/C vdd NAND3X1
XNAND2X1_49 NAND2X1_49/A NAND2X1_49/B gnd OR2X2_8/A vdd NAND2X1
XNAND2X1_38 INVX2_15/Y XOR2X1_4/Y gnd NAND2X1_38/Y vdd NAND2X1
XNAND2X1_27 AND2X2_6/B AND2X2_6/A gnd AND2X2_7/A vdd NAND2X1
XNAND2X1_16 BUFX4_1/Y a[7] gnd NAND3X1_5/C vdd NAND2X1
XAOI22X1_6 BUFX4_1/Y a[4] a[3] BUFX4_14/Y gnd OAI22X1_8/C vdd AOI22X1
XNOR3X1_4 NOR3X1_4/A NOR3X1_4/B NOR3X1_4/C gnd NOR3X1_4/Y vdd NOR3X1
XOAI22X1_9 INVX4_7/Y INVX1_41/Y INVX4_5/Y NOR2X1_64/A gnd OR2X2_10/A vdd OAI22X1
XINVX2_18 INVX2_18/A gnd NOR2X1_3/A vdd INVX2
XXOR2X1_1 XOR2X1_1/A NOR2X1_9/Y gnd XOR2X1_1/Y vdd XOR2X1
XFILL_6_0_0 gnd vdd FILL
XMUX2X1_2 a[3] a[2] BUFX4_3/Y gnd MUX2X1_2/Y vdd MUX2X1
XBUFX4_14 b[1] gnd BUFX4_14/Y vdd BUFX4
XNAND3X1_2 INVX1_4/Y INVX1_5/A OR2X2_1/Y gnd AND2X2_4/B vdd NAND3X1
XAOI22X1_7 INVX1_11/Y INVX2_13/Y AOI22X1_7/C AOI22X1_7/D gnd DFFSR_5/D vdd AOI22X1
XNAND2X1_28 BUFX4_3/Y INVX4_4/Y gnd AND2X2_7/B vdd NAND2X1
XFILL_1_1_1 gnd vdd FILL
XOAI21X1_120 AOI21X1_68/Y AOI21X1_69/Y INVX1_43/Y gnd NAND3X1_66/C vdd OAI21X1
XNAND2X1_17 BUFX4_5/Y a[1] gnd OAI21X1_54/A vdd NAND2X1
XNAND2X1_39 a[3] INVX8_2/A gnd OAI22X1_6/B vdd NAND2X1
XNOR3X1_5 INVX1_32/A INVX1_34/A NOR3X1_5/C gnd NOR3X1_5/Y vdd NOR3X1
XAOI21X1_70 INVX2_20/Y AOI21X1_70/B NOR2X1_61/Y gnd AOI21X1_70/Y vdd AOI21X1
XINVX2_19 INVX2_19/A gnd INVX2_19/Y vdd INVX2
XXOR2X1_2 INVX1_6/A NOR2X1_9/Y gnd XOR2X1_2/Y vdd XOR2X1
XMUX2X1_3 a[4] a[3] BUFX4_5/Y gnd MUX2X1_5/A vdd MUX2X1
XFILL_6_0_1 gnd vdd FILL
XOAI21X1_110 INVX2_23/Y OR2X2_4/Y en gnd OR2X2_10/B vdd OAI21X1
XNAND3X1_3 a[4] b[3] OAI22X1_3/B gnd AND2X2_3/A vdd NAND3X1
XOAI21X1_121 NOR2X1_71/Y OAI22X1_4/C INVX1_43/A gnd NAND3X1_66/B vdd OAI21X1
XAOI22X1_8 BUFX4_3/Y a[5] BUFX4_11/Y a[4] gnd AOI22X1_8/Y vdd AOI22X1
XNOR3X1_6 NOR3X1_6/A OR2X2_8/Y NOR3X1_6/C gnd NOR3X1_6/Y vdd NOR3X1
XNAND2X1_29 INVX4_1/A a[2] gnd INVX2_12/A vdd NAND2X1
XNAND2X1_18 a[0] BUFX4_1/Y gnd INVX2_6/A vdd NAND2X1
XAOI21X1_60 NAND3X1_56/Y NAND3X1_57/C INVX2_19/A gnd NOR3X1_6/A vdd AOI21X1
XAOI21X1_71 NAND3X1_46/B NAND3X1_46/C INVX2_21/Y gnd AOI21X1_72/C vdd AOI21X1
XMUX2X1_4 a[6] a[5] BUFX4_1/Y gnd MUX2X1_5/B vdd MUX2X1
XXOR2X1_3 XOR2X1_3/A OR2X2_1/A gnd XOR2X1_3/Y vdd XOR2X1
XFILL_12_0_0 gnd vdd FILL
XINVX4_1 INVX4_1/A gnd INVX4_1/Y vdd INVX4
XBUFX4_1 b[0] gnd BUFX4_1/Y vdd BUFX4
XFILL_4_1_0 gnd vdd FILL
XAOI22X1_9 INVX1_10/Y INVX2_13/Y NOR2X1_67/Y AOI22X1_9/D gnd DFFSR_6/D vdd AOI22X1
XOAI21X1_100 AOI21X1_54/Y OAI21X1_95/B INVX1_38/Y gnd NAND2X1_58/B vdd OAI21X1
XOAI21X1_122 AOI21X1_66/Y AOI21X1_67/Y INVX1_42/Y gnd NAND2X1_68/A vdd OAI21X1
XNAND3X1_4 a[3] b[4] NAND3X1_4/C gnd AND2X2_3/B vdd NAND3X1
XOAI21X1_111 NOR2X1_66/Y OAI21X1_111/B AOI21X1_64/Y gnd OR2X2_11/B vdd OAI21X1
XNAND2X1_19 opcode[0] INVX1_17/Y gnd NOR2X1_29/B vdd NAND2X1
XAOI21X1_61 NAND3X1_60/Y AOI21X1_61/B INVX2_19/Y gnd NOR3X1_6/C vdd AOI21X1
XFILL_9_0_0 gnd vdd FILL
XAOI21X1_72 NAND3X1_48/A NAND3X1_51/Y AOI21X1_72/C gnd AOI21X1_72/Y vdd AOI21X1
XOAI21X1_1 INVX2_22/Y b[5] OAI21X1_1/C gnd INVX1_1/A vdd OAI21X1
XAOI21X1_50 INVX2_18/A INVX1_35/Y INVX2_7/Y gnd AOI21X1_52/B vdd AOI21X1
XXOR2X1_4 AND2X2_9/A AND2X2_9/B gnd XOR2X1_4/Y vdd XOR2X1
XMUX2X1_5 MUX2X1_5/A MUX2X1_5/B INVX8_2/Y gnd MUX2X1_5/Y vdd MUX2X1
XBUFX4_2 b[0] gnd BUFX4_2/Y vdd BUFX4
XFILL_4_1_1 gnd vdd FILL
XFILL_12_0_1 gnd vdd FILL
XINVX4_2 a[4] gnd INVX4_2/Y vdd INVX4
XOAI21X1_112 AOI21X1_59/Y INVX2_19/Y NAND3X1_57/C gnd NAND3X1_78/B vdd OAI21X1
XOAI21X1_101 OAI21X1_82/A INVX1_33/A NAND3X1_38/Y gnd NAND3X1_59/C vdd OAI21X1
XNAND3X1_5 INVX8_2/A a[6] NAND3X1_5/C gnd NAND3X1_5/Y vdd NAND3X1
XOAI21X1_123 AND2X2_13/Y NOR2X1_70/Y INVX1_42/A gnd NAND2X1_68/B vdd OAI21X1
XFILL_9_0_1 gnd vdd FILL
XOAI21X1_2 INVX1_41/A NOR2X1_64/A NOR2X1_3/A gnd OAI21X1_3/B vdd OAI21X1
XAOI21X1_62 NAND2X1_59/Y OR2X2_9/Y INVX2_7/Y gnd NOR2X1_67/A vdd AOI21X1
XAOI21X1_73 NAND3X1_69/B NAND3X1_69/C AOI21X1_70/Y gnd AOI21X1_9/C vdd AOI21X1
XAOI21X1_51 INVX4_1/A INVX1_16/Y INVX2_9/Y gnd OAI21X1_92/C vdd AOI21X1
XAOI21X1_40 INVX1_24/A AOI21X1_40/B OAI21X1_74/Y gnd AOI21X1_40/Y vdd AOI21X1
XXOR2X1_5 XOR2X1_5/A XOR2X1_5/B gnd XOR2X1_5/Y vdd XOR2X1
XBUFX4_3 b[0] gnd BUFX4_3/Y vdd BUFX4
XINVX4_3 INVX4_3/A gnd INVX4_3/Y vdd INVX4
XNAND3X1_6 BUFX4_2/Y a[7] NAND2X1_7/Y gnd NAND3X1_6/Y vdd NAND3X1
XOAI21X1_102 AOI21X1_59/Y AOI21X1_58/Y INVX2_19/Y gnd NAND3X1_58/C vdd OAI21X1
XOAI21X1_113 NOR2X1_60/B AND2X2_13/B NAND2X1_58/B gnd XOR2X1_5/A vdd OAI21X1
XOAI21X1_124 AOI21X1_9/C AOI21X1_74/Y OAI21X1_18/B gnd NAND3X1_73/C vdd OAI21X1
XAOI21X1_41 INVX2_7/A XNOR2X1_7/Y OR2X2_7/Y gnd AOI22X1_5/C vdd AOI21X1
XAOI21X1_30 a[1] INVX8_2/Y AND2X2_7/Y gnd NOR2X1_50/B vdd AOI21X1
XAOI21X1_52 AOI21X1_52/A AOI21X1_52/B AOI21X1_52/C gnd AOI22X1_7/C vdd AOI21X1
XOAI21X1_3 INVX1_35/Y OAI21X1_3/B INVX1_1/Y gnd OAI21X1_3/Y vdd OAI21X1
XAOI21X1_63 AOI21X1_63/A NAND2X1_60/Y INVX2_8/Y gnd OR2X2_11/A vdd AOI21X1
XAOI21X1_74 NAND3X1_66/B NAND3X1_66/C OAI22X1_10/Y gnd AOI21X1_74/Y vdd AOI21X1
XFILL_10_1_0 gnd vdd FILL
XFILL_7_1_0 gnd vdd FILL
XBUFX4_4 b[0] gnd BUFX4_4/Y vdd BUFX4
XINVX4_4 a[0] gnd INVX4_4/Y vdd INVX4
XNAND3X1_7 INVX1_7/Y NAND3X1_5/Y NAND3X1_6/Y gnd NAND3X1_7/Y vdd NAND3X1
XOAI21X1_103 NOR3X1_6/A NOR3X1_6/C NOR3X1_5/C gnd NAND3X1_61/B vdd OAI21X1
XBUFX2_1 DFFSR_1/Q gnd out[0] vdd BUFX2
XOAI21X1_114 AOI21X1_65/Y NAND3X1_54/A NAND3X1_52/B gnd NAND3X1_71/C vdd OAI21X1
XOAI21X1_125 OAI21X1_20/A AOI21X1_4/C INVX2_25/Y gnd NAND3X1_81/C vdd OAI21X1
XINVX2_1 INVX2_1/A gnd INVX2_1/Y vdd INVX2
XAOI21X1_1 INVX2_9/A AOI21X1_1/B OAI21X1_9/Y gnd AOI21X1_1/Y vdd AOI21X1
XAOI21X1_42 INVX2_14/Y NAND3X1_33/Y AOI21X1_35/Y gnd OR2X2_8/B vdd AOI21X1
XAOI21X1_53 INVX1_33/Y AOI21X1_53/B AOI21X1_53/C gnd AOI21X1_53/Y vdd AOI21X1
XAOI21X1_75 INVX2_19/A NAND3X1_56/Y AOI21X1_58/Y gnd AOI21X1_75/Y vdd AOI21X1
XAOI21X1_31 NOR2X1_50/A NOR2X1_50/B AOI21X1_31/C gnd NOR2X1_45/A vdd AOI21X1
XOAI21X1_4 INVX1_37/Y NOR2X1_64/A INVX1_41/Y gnd NOR2X1_4/A vdd OAI21X1
XAOI21X1_20 OR2X2_2/B OAI21X1_26/A AOI21X1_20/C gnd NOR3X1_4/C vdd AOI21X1
XAOI21X1_64 NAND2X1_24/B INVX1_2/A OR2X2_10/Y gnd AOI21X1_64/Y vdd AOI21X1
XFILL_3_1 gnd vdd FILL
XFILL_10_1_1 gnd vdd FILL
XFILL_7_1_1 gnd vdd FILL
XBUFX4_5 b[0] gnd BUFX4_5/Y vdd BUFX4
XINVX4_5 INVX4_5/A gnd INVX4_5/Y vdd INVX4
XOAI21X1_126 AOI22X1_11/Y AOI21X1_78/Y NAND3X1_64/B gnd NAND3X1_86/B vdd OAI21X1
XOAI21X1_104 NOR3X1_6/A NOR3X1_6/C OR2X2_8/Y gnd NAND3X1_63/C vdd OAI21X1
XBUFX2_2 BUFX2_2/A gnd out[1] vdd BUFX2
XOAI21X1_115 AND2X2_13/Y NOR2X1_70/Y INVX1_42/Y gnd NAND2X1_64/B vdd OAI21X1
XNAND3X1_8 NAND3X1_7/Y AOI21X1_8/B INVX1_6/Y gnd NAND3X1_8/Y vdd NAND3X1
XINVX2_2 INVX2_2/A gnd INVX2_2/Y vdd INVX2
XAOI21X1_2 INVX2_7/A XNOR2X1_1/Y AOI21X1_2/C gnd AOI21X1_2/Y vdd AOI21X1
XAOI21X1_43 INVX2_15/Y OAI21X1_77/Y NOR2X1_48/Y gnd AOI21X1_43/Y vdd AOI21X1
XAOI21X1_54 a[2] b[3] OAI21X1_76/B gnd AOI21X1_54/Y vdd AOI21X1
XAOI21X1_65 NAND3X1_47/A NAND3X1_47/B INVX2_21/A gnd AOI21X1_65/Y vdd AOI21X1
XAOI21X1_76 NAND3X1_71/A NAND3X1_71/B AOI21X1_72/Y gnd AOI21X1_4/C vdd AOI21X1
XOAI21X1_5 NOR2X1_4/Y INVX2_1/Y INVX2_8/A gnd OAI21X1_5/Y vdd OAI21X1
XAOI21X1_10 NAND3X1_7/Y AOI21X1_8/B XOR2X1_1/A gnd OAI21X1_17/B vdd AOI21X1
XAOI21X1_21 OAI21X1_28/Y OR2X2_2/Y INVX2_8/Y gnd NOR3X1_4/A vdd AOI21X1
XAOI21X1_32 BUFX4_6/Y OAI21X1_9/B INVX4_3/Y gnd AOI21X1_32/Y vdd AOI21X1
XINVX4_6 a[2] gnd INVX4_6/Y vdd INVX4
XBUFX4_6 b[2] gnd BUFX4_6/Y vdd BUFX4
XBUFX2_3 BUFX2_3/A gnd out[2] vdd BUFX2
XOAI21X1_116 AOI21X1_66/Y AOI21X1_67/Y INVX1_42/A gnd NAND2X1_64/A vdd OAI21X1
XNAND3X1_9 NAND3X1_8/Y NAND3X1_9/B XNOR2X1_2/Y gnd NAND3X1_9/Y vdd NAND3X1
XOAI21X1_105 INVX4_2/Y b[4] AOI21X1_52/A gnd OR2X2_9/A vdd OAI21X1
XAOI21X1_3 AOI21X1_2/Y AOI21X1_3/B AOI21X1_3/C gnd DFFSR_7/D vdd AOI21X1
XINVX2_3 INVX2_3/A gnd OR2X2_2/B vdd INVX2
XNOR2X1_1 a[6] b[6] gnd NOR2X1_2/A vdd NOR2X1
XAOI21X1_33 INVX1_25/A AOI21X1_33/B NOR2X1_47/Y gnd INVX1_27/A vdd AOI21X1
XAOI21X1_55 a[1] b[4] OAI22X1_3/A gnd OAI21X1_95/B vdd AOI21X1
XAOI21X1_77 NAND3X1_73/A NAND3X1_73/C NAND3X1_71/C gnd OAI21X1_20/A vdd AOI21X1
XAOI21X1_11 NAND3X1_13/A NAND3X1_13/C OAI21X1_18/Y gnd OAI21X1_19/A vdd AOI21X1
XOAI21X1_6 INVX2_4/Y BUFX4_1/Y NOR2X1_61/A gnd NOR2X1_5/B vdd OAI21X1
XAOI21X1_22 NOR2X1_5/A NAND2X1_61/B OAI21X1_29/Y gnd NOR2X1_14/B vdd AOI21X1
XAOI21X1_66 a[3] b[3] AND2X2_13/B gnd AOI21X1_66/Y vdd AOI21X1
XAOI21X1_44 BUFX4_4/Y a[4] OAI22X1_6/B gnd AOI21X1_44/Y vdd AOI21X1
XFILL_2_0_0 gnd vdd FILL
XFILL_13_1 gnd vdd FILL
XBUFX4_7 b[2] gnd BUFX4_7/Y vdd BUFX4
XINVX4_7 INVX4_7/A gnd INVX4_7/Y vdd INVX4
XOAI21X1_106 NOR2X1_65/B INVX1_37/A INVX2_23/Y gnd AOI21X1_63/A vdd OAI21X1
XOAI21X1_117 NOR2X1_71/Y OAI22X1_4/C INVX1_43/Y gnd NAND3X1_69/B vdd OAI21X1
XBUFX2_4 BUFX2_4/A gnd out[3] vdd BUFX2
XAOI21X1_4 XOR2X1_5/Y AOI21X1_4/B AOI21X1_4/C gnd AOI21X1_4/Y vdd AOI21X1
XINVX2_4 a[6] gnd INVX2_4/Y vdd INVX2
XNOR2X1_2 NOR2X1_2/A INVX1_3/A gnd INVX2_1/A vdd NOR2X1
XAOI21X1_78 NAND3X1_78/Y AOI21X1_78/B NAND3X1_63/B gnd AOI21X1_78/Y vdd AOI21X1
XAOI21X1_34 NAND3X1_34/B NAND3X1_33/Y INVX2_14/Y gnd OAI21X1_69/B vdd AOI21X1
XAOI21X1_23 NOR3X1_4/Y NAND3X1_24/Y NOR2X1_17/Y gnd DFFSR_8/D vdd AOI21X1
XAOI21X1_67 a[2] b[4] NOR2X1_70/A gnd AOI21X1_67/Y vdd AOI21X1
XAOI21X1_12 NAND3X1_9/Y NAND3X1_10/C XOR2X1_3/A gnd OAI21X1_19/B vdd AOI21X1
XOAI21X1_7 OAI21X1_7/A INVX8_2/Y INVX4_1/Y gnd OAI21X1_7/Y vdd OAI21X1
XAOI21X1_56 BUFX4_4/Y a[5] OAI22X1_8/B gnd OAI21X1_97/A vdd AOI21X1
XAOI21X1_45 a[3] BUFX4_13/Y NOR2X1_52/A gnd OAI21X1_80/B vdd AOI21X1
XFILL_1_1 gnd vdd FILL
XFILL_2_0_1 gnd vdd FILL
XBUFX4_8 b[2] gnd INVX4_1/A vdd BUFX4
XBUFX2_5 DFFSR_5/Q gnd out[4] vdd BUFX2
XOAI21X1_107 INVX2_22/Y BUFX4_5/Y NOR2X1_52/A gnd NAND2X1_61/B vdd OAI21X1
XOAI21X1_118 AOI21X1_68/Y AOI21X1_69/Y INVX1_43/A gnd NAND3X1_69/C vdd OAI21X1
XINVX2_5 opcode[2] gnd INVX2_5/Y vdd INVX2
XAOI21X1_5 BUFX4_3/Y a[7] NAND2X1_7/Y gnd NOR3X1_1/A vdd AOI21X1
XAOI21X1_35 NAND3X1_33/B OAI21X1_68/Y INVX1_27/A gnd AOI21X1_35/Y vdd AOI21X1
XAOI21X1_46 AOI21X1_46/A AOI21X1_46/B AOI21X1_43/Y gnd AOI21X1_53/C vdd AOI21X1
XNOR2X1_3 NOR2X1_3/A INVX2_23/Y gnd AND2X2_1/B vdd NOR2X1
XAOI21X1_68 BUFX4_3/Y a[6] NOR2X1_71/B gnd AOI21X1_68/Y vdd AOI21X1
XAOI21X1_57 INVX8_2/A a[4] NOR2X1_61/A gnd OAI21X1_97/B vdd AOI21X1
XAOI21X1_24 INVX1_16/A INVX1_24/A OAI21X1_38/Y gnd NAND2X1_21/B vdd AOI21X1
XAOI21X1_13 NAND3X1_19/B NAND3X1_19/C AOI21X1_4/Y gnd NOR2X1_10/A vdd AOI21X1
XAOI21X1_79 NAND3X1_61/A NAND3X1_61/B NAND3X1_42/C gnd AOI21X1_79/Y vdd AOI21X1
XOAI21X1_8 INVX4_7/Y INVX1_3/Y en gnd NOR2X1_6/A vdd OAI21X1
XOAI22X1_10 NOR2X1_52/A NOR2X1_71/B AOI22X1_8/Y INVX2_20/A gnd OAI22X1_10/Y vdd OAI22X1
XFILL_1_2 gnd vdd FILL
XBUFX4_9 b[2] gnd BUFX4_9/Y vdd BUFX4
XBUFX2_6 BUFX2_6/A gnd out[5] vdd BUFX2
XNAND2X1_1 a[0] b[7] gnd INVX1_4/A vdd NAND2X1
XOAI21X1_108 INVX1_40/Y INVX8_2/Y NAND2X1_61/Y gnd NOR2X1_66/B vdd OAI21X1
XOAI21X1_119 INVX8_2/Y INVX4_2/Y NOR2X1_61/A gnd AOI21X1_70/B vdd OAI21X1
XINVX2_6 INVX2_6/A gnd INVX2_6/Y vdd INVX2
XFILL_0_1_0 gnd vdd FILL
XAOI21X1_6 BUFX4_13/Y a[6] NAND3X1_5/C gnd NOR3X1_1/C vdd AOI21X1
XNOR2X1_4 NOR2X1_4/A NOR2X1_4/B gnd NOR2X1_4/Y vdd NOR2X1
XAOI21X1_36 OAI21X1_66/Y NAND2X1_38/Y INVX1_27/Y gnd OAI21X1_70/B vdd AOI21X1
XAOI21X1_58 NAND3X1_48/Y NAND3X1_59/B AOI21X1_53/Y gnd AOI21X1_58/Y vdd AOI21X1
XAOI21X1_47 NAND3X1_38/B NAND3X1_38/A OAI22X1_6/Y gnd OAI21X1_82/A vdd AOI21X1
XAOI21X1_14 NAND3X1_9/Y NAND3X1_10/C INVX1_8/Y gnd AOI21X1_14/Y vdd AOI21X1
XOAI21X1_9 INVX1_2/Y OAI21X1_9/B NOR2X1_6/Y gnd OAI21X1_9/Y vdd OAI21X1
XAOI21X1_69 NOR2X1_5/A a[5] NOR2X1_71/A gnd AOI21X1_69/Y vdd AOI21X1
XAOI21X1_25 NOR2X1_28/Y NAND3X1_29/Y AOI21X1_25/C gnd AOI21X1_25/Y vdd AOI21X1
XFILL_5_0_0 gnd vdd FILL
XBUFX2_7 BUFX2_7/A gnd out[6] vdd BUFX2
XNAND3X1_80 AOI21X1_75/Y NAND3X1_81/B NAND3X1_81/C gnd AOI21X1_78/B vdd NAND3X1
XFILL_11_1 gnd vdd FILL
XOAI21X1_109 AOI22X1_2/B INVX4_1/Y INVX2_9/A gnd OAI21X1_111/B vdd OAI21X1
XFILL_0_1_1 gnd vdd FILL
XAOI21X1_7 NAND3X1_5/Y NAND3X1_6/Y INVX1_7/Y gnd NOR3X1_3/B vdd AOI21X1
XNAND2X1_2 a[3] b[4] gnd OAI22X1_3/B vdd NAND2X1
XINVX2_7 INVX2_7/A gnd INVX2_7/Y vdd INVX2
XNOR2X1_5 NOR2X1_5/A NOR2X1_5/B gnd NOR2X1_5/Y vdd NOR2X1
XAOI21X1_48 NAND2X1_49/B NAND2X1_49/A AOI21X1_48/C gnd INVX1_34/A vdd AOI21X1
XAOI21X1_59 NAND3X1_53/Y NAND3X1_54/Y NAND3X1_59/C gnd AOI21X1_59/Y vdd AOI21X1
XAOI21X1_26 OAI21X1_36/Y AOI21X1_25/Y NOR2X1_21/Y gnd DFFSR_1/D vdd AOI21X1
XAOI21X1_37 NOR2X1_50/A OAI21X1_50/Y INVX2_12/Y gnd INVX1_30/A vdd AOI21X1
XAOI21X1_15 NAND3X1_13/A NAND3X1_13/C INVX1_8/A gnd AOI21X1_15/Y vdd AOI21X1
XFILL_5_0_1 gnd vdd FILL
XBUFX2_8 BUFX2_8/A gnd out[7] vdd BUFX2
XNAND3X1_81 NAND3X1_78/B NAND3X1_81/B NAND3X1_81/C gnd NOR2X1_11/B vdd NAND3X1
XFILL_11_2 gnd vdd FILL
XNAND3X1_70 OAI21X1_18/B NAND3X1_68/Y AOI21X1_9/B gnd NAND3X1_71/B vdd NAND3X1
XNOR2X1_70 NOR2X1_70/A AND2X2_13/B gnd NOR2X1_70/Y vdd NOR2X1
XAOI21X1_8 NAND3X1_7/Y AOI21X1_8/B INVX1_6/Y gnd AOI21X1_8/Y vdd AOI21X1
XINVX2_8 INVX2_8/A gnd INVX2_8/Y vdd INVX2
XNAND2X1_3 OR2X2_1/B OR2X2_1/A gnd INVX1_5/A vdd NAND2X1
XNOR2X1_6 NOR2X1_6/A NOR2X1_6/B gnd NOR2X1_6/Y vdd NOR2X1
XINVX1_40 INVX1_40/A gnd INVX1_40/Y vdd INVX1
XAOI21X1_49 OR2X2_6/B INVX2_16/A NOR2X1_56/Y gnd OAI21X1_86/C vdd AOI21X1
XAOI21X1_27 NOR2X1_5/A MUX2X1_5/A BUFX4_6/Y gnd AOI21X1_27/Y vdd AOI21X1
XAOI21X1_16 NAND3X1_18/B NAND3X1_18/C OAI21X1_20/Y gnd NOR2X1_10/B vdd AOI21X1
XAOI21X1_38 AOI21X1_38/A AOI21X1_38/B INVX2_8/Y gnd OR2X2_7/A vdd AOI21X1
XOAI21X1_90 INVX4_2/Y BUFX4_2/Y AND2X2_9/A gnd OAI21X1_7/A vdd OAI21X1
XFILL_3_1_0 gnd vdd FILL
XFILL_11_0_0 gnd vdd FILL
XNAND3X1_82 NAND3X1_82/A AOI21X1_75/Y NAND3X1_77/Y gnd AOI22X1_11/D vdd NAND3X1
XFILL_11_3 gnd vdd FILL
XNAND3X1_60 NAND3X1_53/Y NAND3X1_54/Y AOI21X1_53/Y gnd NAND3X1_60/Y vdd NAND3X1
XNOR2X1_60 NOR2X1_60/A NOR2X1_60/B gnd INVX2_19/A vdd NOR2X1
XNAND3X1_71 NAND3X1_71/A NAND3X1_71/B NAND3X1_71/C gnd NAND3X1_74/B vdd NAND3X1
XNOR2X1_71 NOR2X1_71/A NOR2X1_71/B gnd NOR2X1_71/Y vdd NOR2X1
XBUFX2_9 BUFX2_9/A gnd zero vdd BUFX2
XINVX2_9 INVX2_9/A gnd INVX2_9/Y vdd INVX2
XNAND2X1_4 AND2X2_4/B AND2X2_4/A gnd NAND2X1_4/Y vdd NAND2X1
XAOI21X1_9 AOI21X1_9/A AOI21X1_9/B AOI21X1_9/C gnd XOR2X1_3/A vdd AOI21X1
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XNOR2X1_7 INVX2_10/Y NOR2X1_7/B gnd OR2X2_1/B vdd NOR2X1
XAOI21X1_17 NAND3X1_78/B NAND2X1_10/Y INVX2_2/A gnd OAI21X1_22/A vdd AOI21X1
XAOI21X1_39 BUFX4_6/Y NOR2X1_15/A INVX4_3/Y gnd AOI21X1_39/Y vdd AOI21X1
XAOI21X1_28 OAI21X1_40/Y NAND2X1_24/Y INVX4_3/Y gnd AOI21X1_28/Y vdd AOI21X1
XFILL_8_0_0 gnd vdd FILL
XOAI21X1_80 AOI21X1_44/Y OAI21X1_80/B INVX2_12/Y gnd NAND3X1_38/A vdd OAI21X1
XOAI21X1_91 INVX1_36/Y INVX8_2/Y OAI21X1_91/C gnd OAI21X1_91/Y vdd OAI21X1
XFILL_3_1_1 gnd vdd FILL
XNAND3X1_61 NAND3X1_61/A NAND3X1_61/B NAND3X1_42/C gnd NAND3X1_61/Y vdd NAND3X1
XNOR2X1_72 NOR3X1_6/A NOR3X1_6/C gnd NOR2X1_72/Y vdd NOR2X1
XNAND3X1_83 NOR2X1_11/B AOI22X1_11/D NOR3X1_6/Y gnd NAND3X1_83/Y vdd NAND3X1
XFILL_11_0_1 gnd vdd FILL
XNOR2X1_50 NOR2X1_50/A NOR2X1_50/B gnd OR2X2_6/A vdd NOR2X1
XNAND3X1_50 INVX2_21/A NAND3X1_47/A NAND3X1_47/B gnd NAND3X1_52/B vdd NAND3X1
XNOR2X1_61 NOR2X1_61/A OAI22X1_8/B gnd NOR2X1_61/Y vdd NOR2X1
XNAND3X1_72 AOI21X1_9/A NAND3X1_68/Y AOI21X1_9/B gnd NAND3X1_73/A vdd NAND3X1
XNAND2X1_5 a[4] b[3] gnd NAND3X1_4/C vdd NAND2X1
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XINVX1_20 BUFX4_2/Y gnd AND2X2_5/A vdd INVX1
XINVX1_31 a[3] gnd INVX1_31/Y vdd INVX1
XAOI21X1_18 NAND3X1_85/B AOI21X1_79/Y AOI21X1_78/Y gnd OAI21X1_23/C vdd AOI21X1
XAOI21X1_29 NOR2X1_50/A OAI21X1_50/Y AOI21X1_29/C gnd OAI21X1_64/B vdd AOI21X1
XNOR2X1_8 OR2X2_1/B OR2X2_1/A gnd NOR2X1_8/Y vdd NOR2X1
XFILL_8_0_1 gnd vdd FILL
XOAI21X1_70 AOI21X1_35/Y OAI21X1_70/B INVX2_14/A gnd OAI21X1_70/Y vdd OAI21X1
XOAI21X1_81 NOR2X1_52/Y OAI22X1_8/C INVX2_12/A gnd NAND3X1_38/B vdd OAI21X1
XOAI21X1_92 OAI21X1_91/Y BUFX4_9/Y OAI21X1_92/C gnd AND2X2_12/B vdd OAI21X1
XNAND3X1_84 NAND3X1_63/B NAND3X1_78/Y AOI21X1_78/B gnd NAND3X1_85/B vdd NAND3X1
XNAND3X1_62 NOR3X1_5/C NAND3X1_58/B NAND3X1_58/C gnd NAND3X1_63/B vdd NAND3X1
XNAND3X1_40 INVX1_33/Y AOI21X1_53/B NAND3X1_38/Y gnd NAND2X1_49/A vdd NAND3X1
XNAND3X1_51 NAND3X1_46/B NAND3X1_46/C INVX2_21/Y gnd NAND3X1_51/Y vdd NAND3X1
XNAND3X1_73 NAND3X1_73/A AOI21X1_72/Y NAND3X1_73/C gnd NAND3X1_73/Y vdd NAND3X1
XNOR2X1_51 BUFX4_9/Y INVX4_6/Y gnd OR2X2_6/B vdd NOR2X1
XNOR2X1_73 INVX2_4/Y NOR2X1_7/B gnd INVX1_3/A vdd NOR2X1
XNOR2X1_62 INVX2_22/Y NOR2X1_9/B gnd INVX1_41/A vdd NOR2X1
XNAND2X1_6 AND2X2_3/A AND2X2_3/B gnd XOR2X1_1/A vdd NAND2X1
XNOR2X1_40 NOR2X1_5/A INVX1_22/Y gnd AOI22X1_2/B vdd NOR2X1
XINVX1_10 BUFX2_6/A gnd INVX1_10/Y vdd INVX1
XINVX1_32 INVX1_32/A gnd INVX1_32/Y vdd INVX1
XINVX1_21 INVX1_21/A gnd INVX1_21/Y vdd INVX1
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XNOR2X1_9 INVX4_6/Y NOR2X1_9/B gnd NOR2X1_9/Y vdd NOR2X1
XAOI21X1_19 NAND2X1_12/Y NAND3X1_20/Y AOI21X1_19/C gnd AOI21X1_19/Y vdd AOI21X1
XOAI21X1_82 OAI21X1_82/A AOI21X1_53/C INVX1_33/A gnd NAND2X1_49/B vdd OAI21X1
XFILL_8_1 gnd vdd FILL
XOAI21X1_93 INVX4_7/Y INVX1_37/Y en gnd NOR2X1_59/A vdd OAI21X1
XOAI21X1_71 MUX2X1_5/Y BUFX4_7/Y AOI21X1_39/Y gnd OAI21X1_71/Y vdd OAI21X1
XOAI21X1_60 MUX2X1_2/Y BUFX4_11/Y NAND2X1_31/Y gnd OAI21X1_60/Y vdd OAI21X1
XFILL_6_1_0 gnd vdd FILL
XNAND3X1_41 OR2X2_8/Y INVX1_34/Y INVX1_32/Y gnd NAND3X1_42/C vdd NAND3X1
XNAND3X1_63 NOR3X1_5/Y NAND3X1_63/B NAND3X1_63/C gnd NAND3X1_64/B vdd NAND3X1
XNAND3X1_85 AOI21X1_79/Y NAND3X1_85/B NAND3X1_83/Y gnd NAND3X1_85/Y vdd NAND3X1
XNAND3X1_52 NAND3X1_54/A NAND3X1_52/B NAND3X1_51/Y gnd NAND3X1_59/B vdd NAND3X1
XNAND3X1_74 XOR2X1_5/Y NAND3X1_74/B NAND3X1_73/Y gnd NAND3X1_82/A vdd NAND3X1
XNOR2X1_52 NOR2X1_52/A OAI22X1_6/B gnd NOR2X1_52/Y vdd NOR2X1
XNOR2X1_63 a[5] b[5] gnd NOR2X1_64/A vdd NOR2X1
XNOR2X1_30 opcode[2] OR2X2_3/Y gnd INVX2_8/A vdd NOR2X1
XNAND2X1_7 BUFX4_11/Y a[6] gnd NAND2X1_7/Y vdd NAND2X1
XNOR2X1_41 BUFX4_9/Y a[2] gnd NOR2X1_42/A vdd NOR2X1
XNAND3X1_30 AOI22X1_3/Y OAI21X1_47/Y AOI22X1_2/Y gnd OR2X2_5/A vdd NAND3X1
XINVX1_11 DFFSR_5/Q gnd INVX1_11/Y vdd INVX1
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XINVX1_22 INVX1_22/A gnd INVX1_22/Y vdd INVX1
XOAI21X1_83 OAI21X1_70/B INVX2_14/A NAND3X1_34/B gnd AOI21X1_48/C vdd OAI21X1
XOAI21X1_50 AND2X2_7/A INVX2_6/A AND2X2_6/B gnd OAI21X1_50/Y vdd OAI21X1
XOAI21X1_94 NOR2X1_65/B OAI21X1_94/B AND2X2_12/Y gnd AOI21X1_52/C vdd OAI21X1
XOAI21X1_61 OAI21X1_60/Y BUFX4_7/Y AOI21X1_32/Y gnd OAI21X1_61/Y vdd OAI21X1
XOAI21X1_72 INVX1_31/Y BUFX4_3/Y NOR2X1_47/B gnd INVX1_40/A vdd OAI21X1
XFILL_6_1_1 gnd vdd FILL
XNAND3X1_42 AND2X2_8/A OAI21X1_84/Y NAND3X1_42/C gnd AOI22X1_7/D vdd NAND3X1
XNAND3X1_64 AND2X2_8/A NAND3X1_64/B NAND3X1_61/Y gnd AOI22X1_9/D vdd NAND3X1
XNAND3X1_86 AND2X2_8/A NAND3X1_86/B NAND3X1_85/Y gnd AOI21X1_3/B vdd NAND3X1
XNOR2X1_53 OR2X2_8/B OR2X2_8/A gnd NOR3X1_5/C vdd NOR2X1
XNOR2X1_20 NOR2X1_20/A NOR2X1_20/B gnd BUFX2_9/A vdd NOR2X1
XNAND3X1_20 NAND3X1_78/B INVX2_2/A NAND2X1_10/Y gnd NAND3X1_20/Y vdd NAND3X1
XNAND3X1_31 AND2X2_8/A NAND3X1_31/B INVX1_26/Y gnd NAND3X1_31/Y vdd NAND3X1
XNAND3X1_53 NAND3X1_48/A NAND3X1_52/B NAND3X1_51/Y gnd NAND3X1_53/Y vdd NAND3X1
XNAND3X1_75 NAND3X1_73/A NAND3X1_71/C NAND3X1_73/C gnd NAND3X1_77/C vdd NAND3X1
XNOR2X1_64 NOR2X1_64/A INVX1_41/A gnd OR2X2_9/B vdd NOR2X1
XNOR2X1_31 opcode[0] INVX1_17/Y gnd INVX1_18/A vdd NOR2X1
XNOR2X1_42 NOR2X1_42/A INVX2_12/Y gnd NOR2X1_50/A vdd NOR2X1
XNAND2X1_8 BUFX4_6/Y a[5] gnd INVX1_7/A vdd NAND2X1
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XINVX1_12 BUFX2_4/A gnd INVX1_12/Y vdd INVX1
XINVX1_23 AND2X2_6/B gnd INVX1_23/Y vdd INVX1
XOAI21X1_84 NOR3X1_5/C INVX1_34/A INVX1_32/A gnd OAI21X1_84/Y vdd OAI21X1
XOAI21X1_51 OAI21X1_50/Y NOR2X1_50/A INVX2_8/A gnd AOI21X1_29/C vdd OAI21X1
XOAI21X1_95 AOI21X1_54/Y OAI21X1_95/B INVX1_38/A gnd NAND2X1_55/B vdd OAI21X1
XOAI21X1_40 BUFX4_11/Y OAI21X1_40/B AOI21X1_27/Y gnd OAI21X1_40/Y vdd OAI21X1
XOAI21X1_73 INVX1_22/Y INVX8_2/Y OAI21X1_73/C gnd AOI21X1_40/B vdd OAI21X1
XOAI21X1_62 INVX4_7/Y INVX2_12/A OAI21X1_61/Y gnd NOR2X1_46/B vdd OAI21X1
XAND2X2_10 AND2X2_1/A INVX2_18/A gnd NOR2X1_65/B vdd AND2X2
XNAND3X1_32 OAI21X1_66/Y INVX1_27/Y NAND2X1_38/Y gnd NAND3X1_34/B vdd NAND3X1
XNOR2X1_21 DFFSR_1/Q en gnd NOR2X1_21/Y vdd NOR2X1
XNAND3X1_54 NAND3X1_54/A NAND3X1_46/Y NAND3X1_48/C gnd NAND3X1_54/Y vdd NAND3X1
XNAND3X1_21 NAND2X1_12/Y NAND3X1_20/Y AOI21X1_19/C gnd NAND3X1_21/Y vdd NAND3X1
XNOR2X1_43 INVX4_4/Y INVX4_1/Y gnd INVX1_25/A vdd NOR2X1
XNAND3X1_76 NAND3X1_71/A NAND3X1_71/B AOI21X1_72/Y gnd AOI21X1_4/B vdd NAND3X1
XNAND3X1_43 a[1] b[4] OAI22X1_3/A gnd NAND3X1_49/B vdd NAND3X1
XNOR2X1_54 INVX4_2/Y INVX2_17/Y gnd INVX1_37/A vdd NOR2X1
XNOR2X1_65 INVX1_37/A NOR2X1_65/B gnd NOR2X1_65/Y vdd NOR2X1
XNAND3X1_10 NAND3X1_9/Y XOR2X1_3/A NAND3X1_10/C gnd NAND3X1_14/A vdd NAND3X1
XNAND3X1_65 OAI22X1_10/Y NAND3X1_69/B NAND3X1_69/C gnd NAND3X1_67/B vdd NAND3X1
XNOR2X1_32 INVX2_5/Y NOR2X1_29/B gnd INVX4_7/A vdd NOR2X1
XNOR2X1_10 NOR2X1_10/A NOR2X1_10/B gnd NOR2X1_10/Y vdd NOR2X1
XNAND2X1_9 XOR2X1_5/B XOR2X1_5/A gnd INVX2_2/A vdd NAND2X1
XINVX1_13 BUFX2_3/A gnd INVX1_13/Y vdd INVX1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XFILL_12_1_0 gnd vdd FILL
XOAI21X1_52 NOR2X1_50/B NOR2X1_50/A INVX2_7/A gnd AOI21X1_31/C vdd OAI21X1
XOAI21X1_41 MUX2X1_5/B BUFX4_13/Y NAND2X1_23/Y gnd NAND2X1_24/B vdd OAI21X1
XOAI21X1_30 NOR2X1_14/Y NOR2X1_15/Y INVX4_1/Y gnd NAND3X1_26/C vdd OAI21X1
XOAI21X1_74 INVX4_7/Y NOR2X1_70/A en gnd OAI21X1_74/Y vdd OAI21X1
XOAI21X1_96 NOR2X1_61/Y AOI22X1_8/Y INVX2_20/Y gnd NAND3X1_46/B vdd OAI21X1
XOAI21X1_85 INVX2_12/Y NOR2X1_42/A INVX2_16/A gnd OAI21X1_86/B vdd OAI21X1
XOAI21X1_63 INVX4_5/Y NOR2X1_42/A OAI21X1_63/C gnd NOR2X1_46/A vdd OAI21X1
XAND2X2_11 NOR2X1_59/Y AND2X2_11/B gnd AND2X2_11/Y vdd AND2X2
XFILL_1_0_0 gnd vdd FILL
XFILL_9_1_0 gnd vdd FILL
XNOR2X1_11 INVX2_2/Y NOR2X1_11/B gnd NOR2X1_11/Y vdd NOR2X1
XNOR2X1_44 INVX1_21/Y NOR2X1_44/B gnd INVX1_26/A vdd NOR2X1
XNAND3X1_33 INVX1_27/A NAND3X1_33/B OAI21X1_68/Y gnd NAND3X1_33/Y vdd NAND3X1
XNAND3X1_55 NAND3X1_53/Y NAND3X1_54/Y NAND3X1_59/C gnd NAND3X1_57/C vdd NAND3X1
XNAND3X1_22 NAND3X1_22/A NAND3X1_21/Y OAI21X1_22/Y gnd NAND3X1_22/Y vdd NAND3X1
XNAND3X1_77 AOI21X1_4/B INVX2_25/Y NAND3X1_77/C gnd NAND3X1_77/Y vdd NAND3X1
XNAND3X1_44 a[2] b[3] OAI21X1_76/B gnd NAND3X1_44/Y vdd NAND3X1
XNOR2X1_55 a[4] b[4] gnd NOR2X1_55/Y vdd NOR2X1
XNAND3X1_11 XOR2X1_1/A NAND3X1_7/Y AOI21X1_8/B gnd NAND3X1_11/Y vdd NAND3X1
XNOR2X1_22 INVX2_5/Y OR2X2_3/Y gnd INVX4_3/A vdd NOR2X1
XNOR2X1_66 INVX4_1/A NOR2X1_66/B gnd NOR2X1_66/Y vdd NOR2X1
XNOR2X1_33 opcode[2] OR2X2_4/A gnd INVX2_9/A vdd NOR2X1
XNAND3X1_66 AOI21X1_70/Y NAND3X1_66/B NAND3X1_66/C gnd NAND3X1_67/C vdd NAND3X1
XINVX1_25 INVX1_25/A gnd INVX1_25/Y vdd INVX1
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XFILL_12_1_1 gnd vdd FILL
XOAI21X1_64 NAND2X1_34/Y OAI21X1_64/B en gnd OAI21X1_64/Y vdd OAI21X1
XOAI21X1_75 INVX4_4/Y INVX2_17/Y NOR2X1_60/B gnd OAI21X1_75/Y vdd OAI21X1
XOAI21X1_42 AND2X2_6/Y INVX2_6/Y INVX2_8/A gnd OAI21X1_44/B vdd OAI21X1
XOAI21X1_53 AND2X2_5/A INVX4_6/Y AND2X2_6/B gnd AOI21X1_33/B vdd OAI21X1
XOAI21X1_20 OAI21X1_20/A INVX2_25/Y NAND3X1_77/C gnd OAI21X1_20/Y vdd OAI21X1
XOAI21X1_31 INVX4_7/Y INVX1_9/A en gnd NOR2X1_16/A vdd OAI21X1
XOAI21X1_97 OAI21X1_97/A OAI21X1_97/B INVX2_20/A gnd NAND3X1_46/C vdd OAI21X1
XOAI21X1_86 NOR2X1_50/B OAI21X1_86/B OAI21X1_86/C gnd INVX1_35/A vdd OAI21X1
XAND2X2_12 AND2X2_11/Y AND2X2_12/B gnd AND2X2_12/Y vdd AND2X2
XFILL_1_0_1 gnd vdd FILL
XFILL_9_1_1 gnd vdd FILL
XNAND3X1_34 INVX2_14/Y NAND3X1_34/B NAND3X1_33/Y gnd INVX1_28/A vdd NAND3X1
XNAND3X1_78 NAND3X1_82/A NAND3X1_78/B NAND3X1_77/Y gnd NAND3X1_78/Y vdd NAND3X1
XNAND3X1_56 NAND3X1_48/Y NAND3X1_59/B AOI21X1_53/Y gnd NAND3X1_56/Y vdd NAND3X1
XNAND3X1_23 NAND3X1_78/B INVX2_2/Y NAND2X1_10/Y gnd AOI22X1_1/D vdd NAND3X1
XNAND3X1_45 INVX1_38/Y NAND3X1_49/B NAND3X1_44/Y gnd NAND3X1_45/Y vdd NAND3X1
XNOR2X1_12 a[7] b[7] gnd OAI22X1_5/D vdd NOR2X1
XNAND3X1_12 XNOR2X1_3/Y NAND3X1_11/Y NAND3X1_12/C gnd NAND3X1_13/A vdd NAND3X1
XNAND3X1_67 AOI21X1_9/A NAND3X1_67/B NAND3X1_67/C gnd NAND3X1_71/A vdd NAND3X1
XNOR2X1_45 NOR2X1_45/A NOR2X1_45/B gnd NOR2X1_45/Y vdd NOR2X1
XNOR2X1_67 NOR2X1_67/A OR2X2_11/Y gnd NOR2X1_67/Y vdd NOR2X1
XNOR2X1_23 BUFX4_4/Y INVX4_4/Y gnd INVX1_15/A vdd NOR2X1
XNOR2X1_34 BUFX4_9/Y INVX2_9/Y gnd INVX1_24/A vdd NOR2X1
XNOR2X1_56 b[3] INVX1_31/Y gnd NOR2X1_56/Y vdd NOR2X1
XINVX1_26 INVX1_26/A gnd INVX1_26/Y vdd INVX1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XOAI21X1_65 INVX1_13/Y en OAI21X1_64/Y gnd DFFSR_3/D vdd OAI21X1
XOAI21X1_76 INVX2_14/A OAI21X1_76/B OAI21X1_75/Y gnd INVX1_33/A vdd OAI21X1
XOAI21X1_54 OAI21X1_54/A AND2X2_9/B AOI21X1_33/B gnd XNOR2X1_6/A vdd OAI21X1
XOAI21X1_43 AND2X2_7/A AND2X2_7/B NOR2X1_37/Y gnd OAI21X1_44/C vdd OAI21X1
XOAI21X1_10 AND2X2_2/Y OAI21X1_5/Y AOI21X1_1/Y gnd AOI21X1_2/C vdd OAI21X1
XOAI21X1_87 INVX1_37/A NOR2X1_55/Y INVX1_35/A gnd AOI21X1_52/A vdd OAI21X1
XOAI21X1_21 AOI21X1_14/Y AOI21X1_15/Y XOR2X1_3/Y gnd NAND3X1_18/B vdd OAI21X1
XOAI21X1_32 INVX4_2/Y BUFX4_5/Y NOR2X1_61/A gnd MUX2X1_1/B vdd OAI21X1
XOAI21X1_98 OAI21X1_97/A OAI21X1_97/B INVX2_20/Y gnd NAND3X1_47/B vdd OAI21X1
XAND2X2_13 NOR2X1_70/A AND2X2_13/B gnd AND2X2_13/Y vdd AND2X2
XNAND3X1_35 INVX1_26/A INVX1_28/A OAI21X1_70/Y gnd INVX1_32/A vdd NAND3X1
XNAND3X1_57 INVX2_19/A NAND3X1_56/Y NAND3X1_57/C gnd NAND3X1_58/B vdd NAND3X1
XNOR2X1_68 BUFX2_7/A en gnd AOI21X1_3/C vdd NOR2X1
XNAND3X1_24 AND2X2_8/A OAI21X1_23/Y NAND3X1_22/Y gnd NAND3X1_24/Y vdd NAND3X1
XNAND3X1_46 INVX2_21/A NAND3X1_46/B NAND3X1_46/C gnd NAND3X1_46/Y vdd NAND3X1
XNAND3X1_79 XOR2X1_5/Y AOI21X1_4/B NAND3X1_77/C gnd NAND3X1_81/B vdd NAND3X1
XNOR2X1_13 OAI22X1_5/D INVX1_9/Y gnd INVX2_3/A vdd NOR2X1
XNOR2X1_57 NOR2X1_55/Y INVX1_37/A gnd INVX2_18/A vdd NOR2X1
XNAND3X1_13 NAND3X1_13/A OAI21X1_18/Y NAND3X1_13/C gnd NAND3X1_13/Y vdd NAND3X1
XNAND3X1_68 OAI22X1_10/Y NAND3X1_66/B NAND3X1_66/C gnd NAND3X1_68/Y vdd NAND3X1
XNOR2X1_24 BUFX4_13/Y INVX1_15/Y gnd INVX1_16/A vdd NOR2X1
XNOR2X1_35 INVX2_5/Y INVX1_18/Y gnd INVX4_5/A vdd NOR2X1
XNOR2X1_46 NOR2X1_46/A NOR2X1_46/B gnd NOR2X1_46/Y vdd NOR2X1
XDFFSR_1 DFFSR_1/Q clk DFFSR_6/R vdd DFFSR_1/D gnd vdd DFFSR
XINVX1_27 INVX1_27/A gnd INVX1_27/Y vdd INVX1
XINVX1_38 INVX1_38/A gnd INVX1_38/Y vdd INVX1
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XOAI21X1_11 AOI22X1_11/Y NAND3X1_64/B NAND3X1_83/Y gnd NAND3X1_22/A vdd OAI21X1
XOAI21X1_22 OAI21X1_22/A NOR2X1_11/Y NOR2X1_10/Y gnd OAI21X1_22/Y vdd OAI21X1
XOAI21X1_55 INVX2_6/A AND2X2_6/B NOR2X1_44/B gnd NAND3X1_31/B vdd OAI21X1
XOAI21X1_66 AND2X2_9/Y NOR2X1_48/Y INVX2_15/A gnd OAI21X1_66/Y vdd OAI21X1
XOAI21X1_44 NOR2X1_36/Y OAI21X1_44/B OAI21X1_44/C gnd OR2X2_5/B vdd OAI21X1
XOAI21X1_77 INVX4_6/Y INVX8_2/Y AND2X2_9/A gnd OAI21X1_77/Y vdd OAI21X1
XOAI21X1_33 INVX2_4/Y BUFX4_2/Y NAND3X1_5/C gnd MUX2X1_1/A vdd OAI21X1
XOAI21X1_99 NOR2X1_61/Y AOI22X1_8/Y INVX2_20/A gnd NAND3X1_47/A vdd OAI21X1
XOAI21X1_88 INVX1_30/A INVX1_29/A NOR2X1_70/A gnd AND2X2_1/A vdd OAI21X1
XFILL_4_0_0 gnd vdd FILL
XFILL_4_1 gnd vdd FILL
XNAND3X1_36 AND2X2_8/A INVX1_32/A OAI21X1_69/Y gnd AOI22X1_5/D vdd NAND3X1
XNAND3X1_58 OR2X2_8/Y NAND3X1_58/B NAND3X1_58/C gnd NAND3X1_61/A vdd NAND3X1
XNOR2X1_47 AND2X2_6/B NOR2X1_47/B gnd NOR2X1_47/Y vdd NOR2X1
XNAND3X1_47 NAND3X1_47/A NAND3X1_47/B INVX2_21/Y gnd NAND3X1_48/C vdd NAND3X1
XNOR2X1_36 INVX2_6/A AND2X2_7/A gnd NOR2X1_36/Y vdd NOR2X1
XNOR2X1_69 INVX4_4/Y NOR2X1_7/B gnd XOR2X1_5/B vdd NOR2X1
XNOR2X1_58 BUFX4_6/Y INVX4_3/Y gnd INVX1_2/A vdd NOR2X1
XNOR2X1_14 INVX2_9/Y NOR2X1_14/B gnd NOR2X1_14/Y vdd NOR2X1
XNAND3X1_14 NAND3X1_14/A NAND2X1_4/Y NAND3X1_13/Y gnd NAND3X1_19/B vdd NAND3X1
XNAND3X1_25 BUFX4_7/Y INVX2_9/A AOI21X1_40/B gnd NAND3X1_26/A vdd NAND3X1
XNAND3X1_69 AOI21X1_70/Y NAND3X1_69/B NAND3X1_69/C gnd AOI21X1_9/B vdd NAND3X1
XNOR2X1_25 NOR2X1_25/A NOR2X1_25/B gnd NOR2X1_25/Y vdd NOR2X1
XDFFSR_2 BUFX2_2/A clk DFFSR_6/R vdd DFFSR_2/D gnd vdd DFFSR
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XINVX1_39 b[5] gnd NOR2X1_9/B vdd INVX1
XINVX1_17 opcode[1] gnd INVX1_17/Y vdd INVX1
XOAI21X1_23 AOI21X1_19/Y AOI22X1_1/Y OAI21X1_23/C gnd OAI21X1_23/Y vdd OAI21X1
XOAI21X1_45 INVX4_4/Y INVX8_2/Y OAI21X1_54/A gnd AND2X2_8/B vdd OAI21X1
XOAI21X1_12 INVX1_5/Y NOR2X1_8/Y INVX1_4/A gnd AND2X2_4/A vdd OAI21X1
XOAI21X1_34 MUX2X1_2/Y INVX8_2/Y INVX1_16/Y gnd NOR2X1_25/B vdd OAI21X1
XOAI21X1_67 AND2X2_9/Y NOR2X1_48/Y INVX2_15/Y gnd NAND3X1_33/B vdd OAI21X1
XOAI21X1_78 AOI21X1_44/Y OAI21X1_80/B INVX2_12/A gnd AOI21X1_46/B vdd OAI21X1
XOAI21X1_89 AND2X2_1/A INVX2_18/A INVX2_8/A gnd OAI21X1_94/B vdd OAI21X1
XOAI21X1_56 INVX4_4/Y BUFX4_5/Y BUFX4_13/Y gnd OAI21X1_56/Y vdd OAI21X1
XFILL_4_0_1 gnd vdd FILL
XFILL_4_2 gnd vdd FILL
XNAND3X1_59 NAND3X1_48/Y NAND3X1_59/B NAND3X1_59/C gnd AOI21X1_61/B vdd NAND3X1
XNOR2X1_48 NOR2X1_47/B OAI22X1_6/B gnd NOR2X1_48/Y vdd NOR2X1
XNAND3X1_48 NAND3X1_48/A NAND3X1_46/Y NAND3X1_48/C gnd NAND3X1_48/Y vdd NAND3X1
XNOR2X1_37 INVX2_7/Y AND2X2_7/Y gnd NOR2X1_37/Y vdd NOR2X1
XNAND3X1_26 NAND3X1_26/A NOR2X1_16/Y NAND3X1_26/C gnd NOR3X1_4/B vdd NAND3X1
XNOR2X1_59 NOR2X1_59/A NOR2X1_59/B gnd NOR2X1_59/Y vdd NOR2X1
XNAND3X1_15 INVX1_8/A NAND3X1_13/A NAND3X1_13/C gnd NAND3X1_15/Y vdd NAND3X1
XNOR2X1_15 NOR2X1_15/A INVX4_3/Y gnd NOR2X1_15/Y vdd NOR2X1
XNOR2X1_26 INVX4_3/Y NOR2X1_25/Y gnd NOR2X1_26/Y vdd NOR2X1
XNAND3X1_37 OAI21X1_71/Y AOI22X1_4/Y AOI21X1_40/Y gnd OR2X2_7/B vdd NAND3X1
XDFFSR_3 BUFX2_3/A clk DFFSR_6/R vdd DFFSR_3/D gnd vdd DFFSR
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XINVX1_29 INVX1_29/A gnd INVX1_29/Y vdd INVX1
XOAI21X1_68 INVX4_1/Y INVX2_10/Y XOR2X1_4/Y gnd OAI21X1_68/Y vdd OAI21X1
XOAI21X1_79 NOR2X1_52/Y OAI22X1_8/C INVX2_12/Y gnd AOI21X1_46/A vdd OAI21X1
XOAI21X1_24 INVX1_3/A NOR2X1_2/A OAI21X1_3/Y gnd OAI21X1_25/C vdd OAI21X1
XOAI21X1_13 NOR3X1_1/A NOR3X1_1/C INVX1_7/A gnd AOI21X1_8/B vdd OAI21X1
XOAI21X1_57 INVX4_6/Y BUFX4_1/Y OAI21X1_54/A gnd INVX1_36/A vdd OAI21X1
XOAI21X1_35 OAI21X1_54/A BUFX4_14/Y INVX4_1/Y gnd NOR2X1_25/A vdd OAI21X1
XOAI21X1_46 INVX2_10/Y BUFX4_4/Y INVX2_6/A gnd INVX1_22/A vdd OAI21X1
XNAND3X1_27 INVX1_10/Y INVX1_11/Y NOR2X1_18/Y gnd NOR2X1_20/A vdd NAND3X1
XNOR2X1_38 INVX2_6/A AND2X2_6/B gnd INVX1_21/A vdd NOR2X1
XNAND3X1_38 NAND3X1_38/A NAND3X1_38/B OAI22X1_6/Y gnd NAND3X1_38/Y vdd NAND3X1
XNAND3X1_49 INVX1_38/A NAND3X1_49/B NAND3X1_44/Y gnd NAND2X1_58/A vdd NAND3X1
XNOR2X1_16 NOR2X1_16/A NOR2X1_16/B gnd NOR2X1_16/Y vdd NOR2X1
XNAND3X1_16 INVX1_8/Y NAND3X1_9/Y NAND3X1_10/C gnd NAND3X1_17/B vdd NAND3X1
XFILL_2_1_0 gnd vdd FILL
XNOR2X1_27 a[0] BUFX4_2/Y gnd NOR2X1_27/Y vdd NOR2X1
XNOR2X1_49 a[3] b[3] gnd INVX1_29/A vdd NOR2X1
XFILL_10_0_0 gnd vdd FILL
XDFFSR_4 BUFX2_4/A clk DFFSR_6/R vdd DFFSR_4/D gnd vdd DFFSR
XINVX1_19 BUFX2_2/A gnd INVX1_19/Y vdd INVX1
XNAND2X1_60 OR2X2_9/B NOR2X1_65/Y gnd NAND2X1_60/Y vdd NAND2X1
XFILL_7_0_0 gnd vdd FILL
XOAI21X1_69 INVX1_28/Y OAI21X1_69/B INVX1_26/Y gnd OAI21X1_69/Y vdd OAI21X1
XOAI21X1_25 INVX2_4/Y b[6] OAI21X1_25/C gnd OAI21X1_26/A vdd OAI21X1
XOAI21X1_14 NOR3X1_1/Y NOR3X1_3/B INVX1_6/A gnd NAND3X1_9/B vdd OAI21X1
XOAI21X1_58 INVX1_36/A BUFX4_14/Y OAI21X1_56/Y gnd OAI22X1_1/A vdd OAI21X1
XOAI21X1_36 INVX4_1/Y INVX1_14/Y NOR2X1_26/Y gnd OAI21X1_36/Y vdd OAI21X1
XOAI21X1_47 a[1] BUFX4_11/Y INVX4_5/A gnd OAI21X1_47/Y vdd OAI21X1
XXNOR2X1_1 OAI21X1_3/Y INVX2_1/A gnd XNOR2X1_1/Y vdd XNOR2X1
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XAND2X2_1 AND2X2_1/A AND2X2_1/B gnd NOR2X1_4/B vdd AND2X2
XFILL_2_1 gnd vdd FILL
XNAND3X1_28 INVX1_12/Y INVX1_13/Y NOR2X1_19/Y gnd NOR2X1_20/B vdd NAND3X1
XNOR2X1_17 BUFX2_8/A en gnd NOR2X1_17/Y vdd NOR2X1
XNAND3X1_39 AOI21X1_43/Y AOI21X1_46/A AOI21X1_46/B gnd AOI21X1_53/B vdd NAND3X1
XNAND3X1_17 NAND3X1_15/Y NAND3X1_17/B XNOR2X1_5/Y gnd NAND3X1_18/C vdd NAND3X1
XNOR2X1_28 NOR2X1_27/Y INVX2_6/Y gnd NOR2X1_28/Y vdd NOR2X1
XFILL_10_0_1 gnd vdd FILL
XFILL_2_1_1 gnd vdd FILL
XNOR2X1_39 opcode[2] INVX1_18/Y gnd AND2X2_8/A vdd NOR2X1
XDFFSR_5 DFFSR_5/Q clk DFFSR_6/R vdd DFFSR_5/D gnd vdd DFFSR
XNAND2X1_61 INVX8_2/Y NAND2X1_61/B gnd NAND2X1_61/Y vdd NAND2X1
XNAND2X1_50 INVX8_2/Y OAI21X1_7/A gnd OAI21X1_91/C vdd NAND2X1
XOAI21X1_59 INVX1_24/Y OAI22X1_1/A NAND3X1_31/Y gnd NOR2X1_45/B vdd OAI21X1
XOAI21X1_48 OR2X2_5/Y AOI21X1_28/Y en gnd OAI21X1_48/Y vdd OAI21X1
XFILL_7_0_1 gnd vdd FILL
XOAI21X1_15 NOR3X1_2/Y AOI21X1_8/Y XOR2X1_1/Y gnd NAND3X1_10/C vdd OAI21X1
XOAI21X1_26 OAI21X1_26/A OR2X2_2/B INVX2_7/A gnd AOI21X1_20/C vdd OAI21X1
XOAI21X1_37 INVX4_7/A INVX1_18/A INVX2_6/Y gnd NAND2X1_21/A vdd OAI21X1
XXNOR2X1_2 XOR2X1_1/A NOR2X1_9/Y gnd XNOR2X1_2/Y vdd XNOR2X1
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XAND2X2_2 NOR2X1_4/Y INVX2_1/Y gnd AND2X2_2/Y vdd AND2X2
XNOR2X1_18 BUFX2_8/A BUFX2_7/A gnd NOR2X1_18/Y vdd NOR2X1
XNOR2X1_29 opcode[2] NOR2X1_29/B gnd INVX2_7/A vdd NOR2X1
XNAND3X1_29 INVX2_8/Y OR2X2_4/Y INVX2_7/Y gnd NAND3X1_29/Y vdd NAND3X1
XNAND3X1_18 OAI21X1_20/Y NAND3X1_18/B NAND3X1_18/C gnd AOI22X1_1/A vdd NAND3X1
XDFFSR_6 BUFX2_6/A clk DFFSR_6/R vdd DFFSR_6/D gnd vdd DFFSR
XNAND2X1_62 a[2] b[4] gnd AND2X2_13/B vdd NAND2X1
XNAND2X1_51 INVX1_14/Y INVX1_2/A gnd AND2X2_11/B vdd NAND2X1
XNAND2X1_40 a[3] b[3] gnd NOR2X1_70/A vdd NAND2X1
XOAI21X1_49 INVX1_19/Y en OAI21X1_48/Y gnd DFFSR_2/D vdd OAI21X1
XOAI21X1_27 NOR2X1_4/Y NOR2X1_2/A INVX1_3/Y gnd OR2X2_2/A vdd OAI21X1
XOAI21X1_16 NOR3X1_1/Y NOR3X1_3/B AND2X2_3/Y gnd NAND3X1_12/C vdd OAI21X1
XOAI21X1_38 INVX4_5/Y NOR2X1_27/Y en gnd OAI21X1_38/Y vdd OAI21X1
XINVX2_20 INVX2_20/A gnd INVX2_20/Y vdd INVX2
XXNOR2X1_3 INVX1_6/A NOR2X1_9/Y gnd XNOR2X1_3/Y vdd XNOR2X1
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XFILL_5_1_0 gnd vdd FILL
XAND2X2_3 AND2X2_3/A AND2X2_3/B gnd AND2X2_3/Y vdd AND2X2
XNOR2X1_19 BUFX2_2/A DFFSR_1/Q gnd NOR2X1_19/Y vdd NOR2X1
XNAND3X1_19 AOI21X1_4/Y NAND3X1_19/B NAND3X1_19/C gnd AOI22X1_1/B vdd NAND3X1
XDFFSR_7 BUFX2_7/A clk DFFSR_6/R vdd DFFSR_7/D gnd vdd DFFSR
XNAND2X1_52 a[0] b[4] gnd NOR2X1_60/A vdd NAND2X1
XNAND2X1_63 a[1] b[5] gnd INVX1_42/A vdd NAND2X1
XNAND2X1_30 a[2] INVX8_2/A gnd AND2X2_9/B vdd NAND2X1
XNAND2X1_41 NOR2X1_70/A INVX1_29/Y gnd INVX2_16/A vdd NAND2X1
XOAI22X1_1 OAI22X1_1/A INVX4_1/Y NOR2X1_5/Y OAI21X1_7/Y gnd AOI21X1_1/B vdd OAI22X1
XINVX2_21 INVX2_21/A gnd INVX2_21/Y vdd INVX2
XINVX2_10 a[1] gnd INVX2_10/Y vdd INVX2
XOAI21X1_28 OAI22X1_5/D INVX1_9/Y OR2X2_2/A gnd OAI21X1_28/Y vdd OAI21X1
XOAI21X1_17 NOR3X1_3/Y OAI21X1_17/B XOR2X1_2/Y gnd NAND3X1_13/C vdd OAI21X1
XOAI21X1_39 INVX2_10/Y BUFX4_4/Y NOR2X1_47/B gnd OAI21X1_40/B vdd OAI21X1
XFILL_12_1 gnd vdd FILL
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XXNOR2X1_4 OR2X2_1/B INVX1_4/A gnd INVX1_8/A vdd XNOR2X1
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XFILL_5_1_1 gnd vdd FILL
XAND2X2_4 AND2X2_4/A AND2X2_4/B gnd AND2X2_4/Y vdd AND2X2
XDFFSR_8 BUFX2_8/A clk DFFSR_6/R vdd DFFSR_8/D gnd vdd DFFSR
XNAND2X1_42 INVX2_16/A INVX1_30/Y gnd AOI21X1_38/B vdd NAND2X1
XNAND2X1_64 NAND2X1_64/A NAND2X1_64/B gnd AOI21X1_9/A vdd NAND2X1
XNAND2X1_31 NOR2X1_5/A MUX2X1_1/B gnd NAND2X1_31/Y vdd NAND2X1
XNAND2X1_20 opcode[1] opcode[0] gnd OR2X2_4/A vdd NAND2X1
XNAND2X1_53 a[0] b[5] gnd INVX1_38/A vdd NAND2X1
XOAI22X1_2 OR2X2_4/Y INVX2_1/Y INVX4_5/Y NOR2X1_2/A gnd NOR2X1_6/B vdd OAI22X1
XINVX2_22 a[5] gnd INVX2_22/Y vdd INVX2
XINVX2_11 OR2X2_4/Y gnd INVX2_11/Y vdd INVX2
XOAI21X1_29 BUFX4_14/Y NOR2X1_71/A NOR2X1_15/A gnd OAI21X1_29/Y vdd OAI21X1
XOAI21X1_18 AOI21X1_74/Y OAI21X1_18/B NAND3X1_68/Y gnd OAI21X1_18/Y vdd OAI21X1
XFILL_12_2 gnd vdd FILL
XOR2X2_10 OR2X2_10/A OR2X2_10/B gnd OR2X2_10/Y vdd OR2X2
XOR2X2_3 opcode[1] opcode[0] gnd OR2X2_3/Y vdd OR2X2
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XXNOR2X1_5 XOR2X1_3/A OR2X2_1/A gnd XNOR2X1_5/Y vdd XNOR2X1
.ends

