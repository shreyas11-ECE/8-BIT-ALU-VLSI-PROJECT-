magic
tech scmos
timestamp 1751429576
<< metal1 >>
rect 1000 1303 1002 1307
rect 1006 1303 1009 1307
rect 1013 1303 1016 1307
rect 70 1272 73 1281
rect 322 1278 337 1281
rect 578 1278 588 1281
rect 1374 1278 1382 1281
rect 54 1268 70 1271
rect 286 1268 313 1271
rect 446 1268 462 1271
rect 606 1268 625 1271
rect 666 1268 673 1271
rect 94 1258 97 1268
rect 622 1262 625 1268
rect 202 1258 209 1261
rect 626 1258 641 1261
rect 950 1258 953 1268
rect 1375 1258 1393 1261
rect 230 1248 238 1251
rect 364 1249 366 1253
rect 746 1248 753 1251
rect 226 1238 241 1241
rect 398 1238 406 1241
rect 238 1228 241 1238
rect 210 1218 211 1222
rect 480 1203 482 1207
rect 486 1203 489 1207
rect 493 1203 496 1207
rect 405 1188 406 1192
rect 549 1188 550 1192
rect 102 1168 126 1171
rect 162 1168 169 1171
rect 274 1168 275 1172
rect 722 1168 723 1172
rect 1021 1168 1022 1172
rect 1114 1168 1129 1171
rect 126 1166 130 1168
rect 102 1162 106 1164
rect 146 1158 153 1161
rect 70 1142 73 1151
rect 198 1148 217 1151
rect 266 1148 273 1151
rect 478 1148 505 1151
rect 526 1148 545 1151
rect 622 1148 633 1151
rect 702 1148 710 1151
rect 794 1148 801 1151
rect 1002 1148 1017 1151
rect 1174 1142 1177 1151
rect 1410 1148 1417 1151
rect 222 1138 230 1141
rect 558 1138 574 1141
rect 602 1138 609 1141
rect 782 1138 793 1141
rect 1046 1138 1054 1141
rect 1383 1138 1390 1141
rect 542 1131 545 1138
rect 530 1128 545 1131
rect 558 1128 561 1138
rect 1102 1118 1110 1121
rect 1000 1103 1002 1107
rect 1006 1103 1009 1107
rect 1013 1103 1016 1107
rect 306 1088 313 1091
rect 434 1088 441 1091
rect 842 1088 849 1091
rect 790 1078 798 1081
rect 934 1078 953 1081
rect 966 1078 977 1081
rect 1398 1078 1417 1081
rect 30 1068 49 1071
rect 246 1071 249 1078
rect 966 1072 969 1078
rect 166 1068 177 1071
rect 236 1068 249 1071
rect 730 1068 737 1071
rect 22 1058 30 1061
rect 286 1058 298 1061
rect 414 1058 426 1061
rect 478 1058 486 1061
rect 554 1058 569 1061
rect 582 1058 590 1061
rect 758 1058 769 1061
rect 1006 1058 1022 1061
rect 1222 1058 1230 1061
rect 1418 1058 1425 1061
rect 1462 1061 1465 1068
rect 1454 1058 1465 1061
rect 254 1056 258 1058
rect 294 1056 298 1058
rect 422 1056 426 1058
rect 98 1048 105 1051
rect 566 1048 569 1058
rect 758 1052 761 1058
rect 830 1048 838 1051
rect 21 1038 22 1042
rect 78 1038 118 1041
rect 549 1038 550 1042
rect 1398 1038 1406 1041
rect 480 1003 482 1007
rect 486 1003 489 1007
rect 493 1003 496 1007
rect 226 988 227 992
rect 829 988 830 992
rect 858 988 859 992
rect 909 988 910 992
rect 1162 988 1163 992
rect 1450 988 1451 992
rect 382 972 385 981
rect 966 972 969 981
rect 446 968 470 971
rect 786 968 787 972
rect 90 958 97 961
rect 102 951 105 961
rect 870 958 881 961
rect 994 958 998 962
rect 1006 958 1022 961
rect 870 952 873 958
rect 102 948 110 951
rect 718 942 721 951
rect 770 948 785 951
rect 834 948 857 951
rect 1126 951 1129 961
rect 1110 948 1129 951
rect 1134 948 1153 951
rect 1410 948 1417 951
rect 198 938 217 941
rect 670 938 678 941
rect 766 938 774 941
rect 842 938 849 941
rect 1054 938 1057 948
rect 1150 938 1153 948
rect 1206 938 1225 941
rect 750 931 753 938
rect 750 928 761 931
rect 766 928 769 938
rect 930 928 937 931
rect 1070 928 1089 931
rect 1206 928 1209 938
rect 1000 903 1002 907
rect 1006 903 1009 907
rect 1013 903 1016 907
rect 437 888 438 892
rect 514 888 515 892
rect 788 888 790 892
rect 1026 888 1028 892
rect 406 878 414 882
rect 614 878 622 882
rect 958 878 977 881
rect 1134 878 1145 881
rect 1178 878 1185 881
rect 406 872 409 878
rect 614 872 617 878
rect 270 862 273 871
rect 378 868 385 871
rect 694 868 702 871
rect 810 868 817 871
rect 910 868 918 871
rect 982 868 1009 871
rect 1170 868 1177 871
rect 1222 868 1230 871
rect 1438 868 1449 871
rect 294 858 302 861
rect 450 858 465 861
rect 470 858 478 861
rect 530 858 537 861
rect 686 858 694 861
rect 698 858 713 861
rect 942 858 961 861
rect 1158 858 1166 861
rect 1174 858 1177 868
rect 1290 858 1302 861
rect 1356 858 1358 862
rect 254 848 257 858
rect 142 838 158 841
rect 325 838 326 842
rect 538 838 539 842
rect 480 803 482 807
rect 486 803 489 807
rect 493 803 496 807
rect 645 788 646 792
rect 674 788 675 792
rect 706 788 707 792
rect 730 788 731 792
rect 877 788 878 792
rect 1189 788 1190 792
rect 1413 788 1414 792
rect 758 768 766 771
rect 1378 768 1379 772
rect 38 752 41 761
rect 202 758 206 762
rect 254 751 257 761
rect 282 758 297 761
rect 338 758 342 762
rect 538 758 545 761
rect 238 748 257 751
rect 310 748 334 751
rect 650 748 673 751
rect 806 748 825 751
rect 830 748 849 751
rect 866 748 873 751
rect 974 748 985 751
rect 1174 751 1177 761
rect 1158 748 1177 751
rect 1206 751 1209 761
rect 1494 758 1502 761
rect 1202 748 1209 751
rect 294 738 297 748
rect 806 742 809 748
rect 830 742 833 748
rect 322 738 329 741
rect 386 738 393 741
rect 654 738 662 741
rect 862 738 870 741
rect 1006 738 1030 741
rect 1090 738 1097 741
rect 1198 738 1217 741
rect 1298 738 1305 741
rect 1310 738 1318 741
rect 1358 738 1361 748
rect 1474 738 1481 741
rect 942 732 945 738
rect 938 728 945 732
rect 1310 728 1313 738
rect 994 718 995 722
rect 1490 718 1491 722
rect 1000 703 1002 707
rect 1006 703 1009 707
rect 1013 703 1016 707
rect 130 688 132 692
rect 170 688 177 691
rect 714 688 715 692
rect 733 688 734 692
rect 1058 688 1059 692
rect 1428 688 1430 692
rect 38 671 41 681
rect 58 678 65 681
rect 286 678 294 682
rect 610 678 614 682
rect 286 672 289 678
rect 22 668 41 671
rect 358 668 366 671
rect 414 668 422 671
rect 478 668 502 671
rect 590 668 598 671
rect 826 668 833 671
rect 910 668 921 671
rect 1154 668 1161 671
rect 1198 668 1214 671
rect 1462 671 1465 681
rect 1462 668 1481 671
rect 54 658 65 661
rect 238 661 241 668
rect 246 661 250 664
rect 238 658 250 661
rect 406 658 430 661
rect 470 658 510 661
rect 754 658 761 661
rect 778 658 785 661
rect 910 658 918 661
rect 1030 658 1046 661
rect 1086 658 1113 661
rect 1130 658 1137 661
rect 1274 658 1281 661
rect 446 648 454 651
rect 722 648 729 651
rect 134 638 166 641
rect 902 641 905 648
rect 170 638 177 641
rect 894 638 905 641
rect 258 628 259 632
rect 762 618 763 622
rect 930 618 931 622
rect 1085 618 1086 622
rect 480 603 482 607
rect 486 603 489 607
rect 493 603 496 607
rect 133 588 134 592
rect 498 588 505 591
rect 562 588 563 592
rect 1170 588 1171 592
rect 789 568 790 572
rect 822 566 826 568
rect 14 558 25 561
rect 118 551 121 561
rect 810 558 817 561
rect 1018 558 1022 562
rect 1030 558 1049 561
rect 102 548 121 551
rect 478 548 505 551
rect 514 548 521 551
rect 710 548 721 551
rect 794 548 809 551
rect 970 548 977 551
rect 1058 548 1065 551
rect 1414 551 1417 561
rect 1394 548 1401 551
rect 1414 548 1433 551
rect 1438 548 1446 551
rect 1466 548 1473 551
rect 406 538 414 541
rect 702 538 713 541
rect 806 538 809 548
rect 886 541 889 548
rect 878 538 889 541
rect 1046 538 1054 541
rect 1386 538 1393 541
rect 1426 538 1433 541
rect 710 532 713 538
rect 426 528 430 532
rect 726 528 745 531
rect 878 528 889 531
rect 958 528 969 531
rect 1134 528 1145 531
rect 1294 528 1305 531
rect 1202 518 1203 522
rect 1000 503 1002 507
rect 1006 503 1009 507
rect 1013 503 1016 507
rect 66 488 68 492
rect 106 488 107 492
rect 106 478 121 481
rect 462 478 470 482
rect 726 478 734 482
rect 1422 478 1438 481
rect 166 471 169 478
rect 462 472 465 478
rect 726 472 729 478
rect 126 468 137 471
rect 166 468 177 471
rect 266 468 281 471
rect 334 468 342 471
rect 434 468 441 471
rect 498 468 513 471
rect 578 468 585 471
rect 630 468 649 471
rect 686 468 702 471
rect 926 468 934 471
rect 54 461 57 468
rect 46 458 57 461
rect 326 458 350 461
rect 666 458 673 461
rect 834 458 846 461
rect 950 461 953 471
rect 1134 468 1153 471
rect 1266 468 1273 471
rect 1390 468 1398 471
rect 1446 468 1457 471
rect 926 458 945 461
rect 950 458 969 461
rect 974 458 998 461
rect 1142 458 1150 461
rect 1218 458 1225 461
rect 1262 458 1270 461
rect 1470 458 1497 461
rect 146 448 150 452
rect 370 448 377 451
rect 746 448 753 451
rect 926 448 929 458
rect 950 452 953 458
rect 982 448 990 451
rect 1318 446 1322 448
rect 70 438 78 441
rect 765 418 766 422
rect 1090 418 1091 422
rect 1162 418 1163 422
rect 480 403 482 407
rect 486 403 489 407
rect 493 403 496 407
rect 21 388 22 392
rect 114 388 115 392
rect 762 388 763 392
rect 1290 388 1291 392
rect 1085 378 1086 382
rect 250 358 255 362
rect 774 358 785 361
rect 198 351 202 354
rect 838 352 841 361
rect 1046 361 1049 368
rect 1038 358 1049 361
rect 166 342 169 351
rect 190 348 202 351
rect 414 341 417 351
rect 518 348 526 351
rect 622 348 633 351
rect 678 348 686 351
rect 934 348 953 351
rect 1006 348 1014 351
rect 1086 348 1094 351
rect 1110 348 1121 351
rect 1162 348 1169 351
rect 1194 348 1201 351
rect 1294 348 1305 351
rect 1442 348 1449 351
rect 398 338 417 341
rect 442 338 454 341
rect 482 338 505 341
rect 542 338 550 341
rect 630 341 633 348
rect 630 338 649 341
rect 722 338 729 341
rect 950 338 953 348
rect 1118 342 1121 348
rect 998 338 1022 341
rect 1238 338 1257 341
rect 1262 338 1281 341
rect 1478 338 1486 341
rect 661 328 662 332
rect 1278 328 1281 338
rect 1406 328 1414 331
rect 1000 303 1002 307
rect 1006 303 1009 307
rect 1013 303 1016 307
rect 741 288 742 292
rect 1494 288 1502 291
rect 122 278 129 281
rect 134 278 145 281
rect 910 278 929 281
rect 134 268 142 271
rect 214 268 222 271
rect 298 268 305 271
rect 354 268 361 271
rect 466 268 473 271
rect 614 268 633 271
rect 894 268 905 271
rect 982 268 998 271
rect 1186 268 1193 271
rect 1250 268 1257 271
rect 1294 268 1302 271
rect 1454 271 1457 278
rect 1434 268 1449 271
rect 1454 268 1473 271
rect 318 258 326 261
rect 486 258 502 261
rect 542 258 561 261
rect 574 258 582 261
rect 666 258 673 261
rect 714 258 729 261
rect 886 258 894 261
rect 1206 258 1233 261
rect 1330 258 1345 261
rect 1350 258 1369 261
rect 1418 258 1425 261
rect 1454 258 1462 261
rect 222 248 225 258
rect 558 248 561 258
rect 658 248 665 251
rect 1058 248 1065 251
rect 1074 248 1078 252
rect 36 238 38 242
rect 70 238 86 241
rect 1302 241 1306 244
rect 1302 238 1313 241
rect 370 218 371 222
rect 773 218 774 222
rect 480 203 482 207
rect 486 203 489 207
rect 493 203 496 207
rect 85 188 86 192
rect 597 188 598 192
rect 149 178 150 182
rect 238 171 241 181
rect 222 168 241 171
rect 746 168 753 171
rect 1058 168 1059 172
rect 1157 168 1158 172
rect 1202 168 1209 171
rect 222 158 225 168
rect 770 158 777 161
rect 734 152 738 154
rect 1102 152 1105 161
rect 1386 158 1391 162
rect 86 148 105 151
rect 150 148 174 151
rect 630 148 638 151
rect 698 148 713 151
rect 838 148 862 151
rect 162 138 169 141
rect 418 138 425 141
rect 446 138 454 141
rect 694 138 702 141
rect 726 138 729 148
rect 910 142 913 151
rect 966 148 977 151
rect 1018 148 1033 151
rect 1038 148 1046 151
rect 1074 148 1089 151
rect 1262 148 1270 151
rect 1290 148 1297 151
rect 1354 148 1361 151
rect 966 138 969 148
rect 1198 138 1206 141
rect 1238 138 1257 141
rect 1266 138 1273 141
rect 1340 138 1350 141
rect 1426 138 1433 141
rect 642 128 649 131
rect 694 128 697 138
rect 934 128 945 131
rect 1222 128 1233 131
rect 1494 128 1502 131
rect 306 118 307 122
rect 1000 103 1002 107
rect 1006 103 1009 107
rect 1013 103 1016 107
rect 82 88 84 92
rect 130 88 143 91
rect 586 88 587 92
rect 110 68 118 71
rect 158 68 174 71
rect 454 71 457 81
rect 686 78 694 81
rect 878 78 889 81
rect 1078 78 1089 81
rect 1266 78 1278 81
rect 454 68 470 71
rect 558 68 566 71
rect 614 68 633 71
rect 862 71 865 78
rect 854 68 865 71
rect 1038 68 1057 71
rect 1198 62 1201 71
rect 1234 68 1241 71
rect 1250 68 1257 71
rect 1318 68 1326 71
rect 1334 68 1353 71
rect 1358 68 1374 71
rect 1390 68 1409 71
rect 438 58 478 61
rect 498 58 529 61
rect 710 58 721 61
rect 738 58 745 61
rect 754 58 769 61
rect 838 58 846 61
rect 906 58 921 61
rect 974 58 990 61
rect 1034 58 1041 61
rect 1122 58 1137 61
rect 1246 58 1254 61
rect 1286 58 1302 61
rect 306 48 311 52
rect 402 48 417 51
rect 494 48 497 58
rect 802 48 806 52
rect 886 48 889 58
rect 918 48 921 58
rect 1486 48 1494 51
rect 518 42 522 44
rect 590 42 594 44
rect 480 3 482 7
rect 486 3 489 7
rect 493 3 496 7
<< m2contact >>
rect 1002 1303 1006 1307
rect 1009 1303 1013 1307
rect 470 1288 474 1292
rect 62 1278 66 1282
rect 318 1278 322 1282
rect 478 1278 482 1282
rect 574 1278 578 1282
rect 614 1278 618 1282
rect 662 1278 666 1282
rect 718 1278 722 1282
rect 910 1278 914 1282
rect 1102 1278 1106 1282
rect 1206 1278 1210 1282
rect 1294 1278 1298 1282
rect 1382 1278 1386 1282
rect 1454 1278 1458 1282
rect 46 1268 50 1272
rect 70 1268 74 1272
rect 86 1268 90 1272
rect 94 1268 98 1272
rect 134 1268 138 1272
rect 158 1268 162 1272
rect 198 1268 202 1272
rect 270 1268 274 1272
rect 278 1268 282 1272
rect 342 1268 346 1272
rect 422 1268 426 1272
rect 462 1268 466 1272
rect 630 1268 634 1272
rect 654 1268 658 1272
rect 662 1268 666 1272
rect 782 1268 786 1272
rect 790 1268 794 1272
rect 894 1268 898 1272
rect 950 1268 954 1272
rect 1086 1268 1090 1272
rect 1278 1268 1282 1272
rect 1430 1268 1434 1272
rect 1462 1268 1466 1272
rect 1494 1268 1498 1272
rect 6 1258 10 1262
rect 22 1258 26 1262
rect 38 1258 42 1262
rect 110 1258 114 1262
rect 142 1258 146 1262
rect 182 1258 186 1262
rect 198 1258 202 1262
rect 238 1258 242 1262
rect 262 1258 266 1262
rect 294 1258 298 1262
rect 302 1258 306 1262
rect 350 1258 354 1262
rect 406 1258 410 1262
rect 430 1258 434 1262
rect 454 1258 458 1262
rect 510 1258 514 1262
rect 550 1258 554 1262
rect 598 1258 602 1262
rect 622 1258 626 1262
rect 686 1258 690 1262
rect 742 1258 746 1262
rect 814 1258 818 1262
rect 846 1258 850 1262
rect 1038 1258 1042 1262
rect 1230 1258 1234 1262
rect 1246 1258 1250 1262
rect 1414 1258 1418 1262
rect 1438 1258 1442 1262
rect 30 1248 34 1252
rect 102 1248 106 1252
rect 126 1248 130 1252
rect 158 1248 162 1252
rect 190 1248 194 1252
rect 238 1248 242 1252
rect 366 1249 370 1253
rect 390 1248 394 1252
rect 414 1248 418 1252
rect 446 1248 450 1252
rect 502 1248 506 1252
rect 558 1248 562 1252
rect 654 1248 658 1252
rect 678 1248 682 1252
rect 710 1248 714 1252
rect 742 1248 746 1252
rect 822 1248 826 1252
rect 862 1250 866 1254
rect 1038 1248 1042 1252
rect 1230 1248 1234 1252
rect 1478 1248 1482 1252
rect 14 1238 18 1242
rect 118 1238 122 1242
rect 174 1238 178 1242
rect 222 1238 226 1242
rect 246 1238 250 1242
rect 406 1238 410 1242
rect 518 1238 522 1242
rect 526 1238 530 1242
rect 542 1238 546 1242
rect 694 1238 698 1242
rect 702 1238 706 1242
rect 734 1238 738 1242
rect 806 1238 810 1242
rect 862 1227 866 1231
rect 1406 1228 1410 1232
rect 70 1218 74 1222
rect 182 1218 186 1222
rect 206 1218 210 1222
rect 550 1218 554 1222
rect 742 1218 746 1222
rect 814 1218 818 1222
rect 990 1218 994 1222
rect 1038 1218 1042 1222
rect 1182 1218 1186 1222
rect 1198 1218 1202 1222
rect 1230 1218 1234 1222
rect 1470 1218 1474 1222
rect 1486 1218 1490 1222
rect 482 1203 486 1207
rect 489 1203 493 1207
rect 22 1188 26 1192
rect 94 1188 98 1192
rect 174 1188 178 1192
rect 318 1188 322 1192
rect 382 1188 386 1192
rect 406 1188 410 1192
rect 446 1188 450 1192
rect 550 1188 554 1192
rect 590 1188 594 1192
rect 646 1188 650 1192
rect 758 1188 762 1192
rect 838 1188 842 1192
rect 1062 1188 1066 1192
rect 1166 1188 1170 1192
rect 1254 1188 1258 1192
rect 1478 1188 1482 1192
rect 1430 1178 1434 1182
rect 14 1168 18 1172
rect 46 1168 50 1172
rect 126 1168 130 1172
rect 158 1168 162 1172
rect 254 1168 258 1172
rect 270 1168 274 1172
rect 334 1168 338 1172
rect 374 1168 378 1172
rect 438 1168 442 1172
rect 694 1168 698 1172
rect 718 1168 722 1172
rect 750 1168 754 1172
rect 1022 1168 1026 1172
rect 1102 1168 1106 1172
rect 1110 1168 1114 1172
rect 30 1158 34 1162
rect 62 1158 66 1162
rect 102 1158 106 1162
rect 118 1158 122 1162
rect 142 1158 146 1162
rect 182 1158 186 1162
rect 286 1158 290 1162
rect 350 1158 354 1162
rect 358 1158 362 1162
rect 390 1158 394 1162
rect 422 1158 426 1162
rect 534 1158 538 1162
rect 678 1158 682 1162
rect 734 1158 738 1162
rect 766 1158 770 1162
rect 814 1158 818 1162
rect 838 1158 842 1162
rect 1118 1158 1122 1162
rect 1206 1158 1210 1162
rect 1254 1156 1258 1160
rect 22 1148 26 1152
rect 38 1148 42 1152
rect 54 1148 58 1152
rect 110 1148 114 1152
rect 166 1148 170 1152
rect 230 1148 234 1152
rect 262 1148 266 1152
rect 294 1148 298 1152
rect 342 1148 346 1152
rect 366 1148 370 1152
rect 406 1148 410 1152
rect 430 1148 434 1152
rect 670 1148 674 1152
rect 686 1148 690 1152
rect 710 1148 714 1152
rect 718 1148 722 1152
rect 758 1148 762 1152
rect 790 1148 794 1152
rect 806 1148 810 1152
rect 846 1148 850 1152
rect 998 1148 1002 1152
rect 1054 1148 1058 1152
rect 1086 1148 1090 1152
rect 1110 1148 1114 1152
rect 1142 1148 1146 1152
rect 1182 1148 1186 1152
rect 1214 1148 1218 1152
rect 1246 1148 1250 1152
rect 1406 1148 1410 1152
rect 1438 1148 1442 1152
rect 1462 1148 1466 1152
rect 70 1138 74 1142
rect 142 1138 146 1142
rect 206 1138 210 1142
rect 214 1138 218 1142
rect 230 1138 234 1142
rect 238 1138 242 1142
rect 262 1138 266 1142
rect 302 1138 306 1142
rect 334 1138 338 1142
rect 414 1138 418 1142
rect 470 1138 474 1142
rect 518 1138 522 1142
rect 542 1138 546 1142
rect 574 1138 578 1142
rect 598 1138 602 1142
rect 614 1138 618 1142
rect 638 1138 642 1142
rect 662 1138 666 1142
rect 710 1138 714 1142
rect 886 1138 890 1142
rect 1038 1138 1042 1142
rect 1054 1138 1058 1142
rect 1062 1138 1066 1142
rect 1078 1138 1082 1142
rect 1150 1138 1154 1142
rect 1166 1138 1170 1142
rect 1174 1138 1178 1142
rect 1190 1138 1194 1142
rect 1206 1138 1210 1142
rect 1286 1138 1290 1142
rect 1390 1138 1394 1142
rect 1454 1138 1458 1142
rect 86 1128 90 1132
rect 182 1128 186 1132
rect 254 1128 258 1132
rect 318 1128 322 1132
rect 454 1128 458 1132
rect 510 1128 514 1132
rect 566 1128 570 1132
rect 598 1128 602 1132
rect 630 1128 634 1132
rect 646 1128 650 1132
rect 774 1128 778 1132
rect 902 1128 906 1132
rect 1030 1128 1034 1132
rect 1134 1128 1138 1132
rect 1302 1128 1306 1132
rect 1406 1128 1410 1132
rect 78 1118 82 1122
rect 126 1118 130 1122
rect 462 1118 466 1122
rect 502 1118 506 1122
rect 982 1118 986 1122
rect 1110 1118 1114 1122
rect 1398 1118 1402 1122
rect 1002 1103 1006 1107
rect 1009 1103 1013 1107
rect 166 1088 170 1092
rect 270 1088 274 1092
rect 302 1088 306 1092
rect 366 1088 370 1092
rect 398 1088 402 1092
rect 430 1088 434 1092
rect 518 1088 522 1092
rect 614 1088 618 1092
rect 662 1088 666 1092
rect 806 1088 810 1092
rect 838 1088 842 1092
rect 870 1088 874 1092
rect 894 1088 898 1092
rect 926 1088 930 1092
rect 998 1088 1002 1092
rect 1470 1088 1474 1092
rect 38 1078 42 1082
rect 246 1078 250 1082
rect 262 1078 266 1082
rect 358 1078 362 1082
rect 390 1078 394 1082
rect 622 1078 626 1082
rect 726 1078 730 1082
rect 782 1078 786 1082
rect 798 1078 802 1082
rect 862 1078 866 1082
rect 902 1078 906 1082
rect 958 1078 962 1082
rect 982 1078 986 1082
rect 990 1078 994 1082
rect 1110 1078 1114 1082
rect 1206 1078 1210 1082
rect 1318 1078 1322 1082
rect 1462 1078 1466 1082
rect 54 1068 58 1072
rect 134 1068 138 1072
rect 158 1068 162 1072
rect 278 1068 282 1072
rect 374 1068 378 1072
rect 406 1068 410 1072
rect 558 1068 562 1072
rect 590 1068 594 1072
rect 606 1068 610 1072
rect 630 1068 634 1072
rect 646 1068 650 1072
rect 686 1068 690 1072
rect 726 1068 730 1072
rect 742 1068 746 1072
rect 758 1068 762 1072
rect 814 1068 818 1072
rect 886 1068 890 1072
rect 918 1068 922 1072
rect 966 1068 970 1072
rect 1094 1068 1098 1072
rect 1230 1068 1234 1072
rect 1302 1068 1306 1072
rect 1462 1068 1466 1072
rect 30 1058 34 1062
rect 62 1058 66 1062
rect 86 1058 90 1062
rect 110 1058 114 1062
rect 214 1058 218 1062
rect 246 1058 250 1062
rect 254 1058 258 1062
rect 302 1058 306 1062
rect 334 1058 338 1062
rect 382 1058 386 1062
rect 430 1058 434 1062
rect 462 1058 466 1062
rect 486 1058 490 1062
rect 510 1058 514 1062
rect 550 1058 554 1062
rect 574 1058 578 1062
rect 590 1058 594 1062
rect 598 1058 602 1062
rect 638 1058 642 1062
rect 678 1058 682 1062
rect 710 1058 714 1062
rect 750 1058 754 1062
rect 822 1058 826 1062
rect 838 1058 842 1062
rect 878 1058 882 1062
rect 910 1058 914 1062
rect 942 1058 946 1062
rect 966 1058 970 1062
rect 1022 1058 1026 1062
rect 1150 1058 1154 1062
rect 1230 1058 1234 1062
rect 1246 1058 1250 1062
rect 1270 1058 1274 1062
rect 1414 1058 1418 1062
rect 1438 1058 1442 1062
rect 1478 1058 1482 1062
rect 6 1048 10 1052
rect 94 1048 98 1052
rect 150 1048 154 1052
rect 190 1048 194 1052
rect 222 1048 226 1052
rect 294 1048 298 1052
rect 326 1048 330 1052
rect 350 1048 354 1052
rect 422 1048 426 1052
rect 454 1048 458 1052
rect 502 1048 506 1052
rect 534 1048 538 1052
rect 654 1048 658 1052
rect 662 1048 666 1052
rect 694 1048 698 1052
rect 718 1048 722 1052
rect 758 1048 762 1052
rect 774 1048 778 1052
rect 838 1048 842 1052
rect 1062 1050 1066 1054
rect 1206 1048 1210 1052
rect 1254 1048 1258 1052
rect 1430 1048 1434 1052
rect 22 1038 26 1042
rect 118 1038 122 1042
rect 206 1038 210 1042
rect 238 1038 242 1042
rect 310 1038 314 1042
rect 342 1038 346 1042
rect 438 1038 442 1042
rect 470 1038 474 1042
rect 518 1038 522 1042
rect 550 1038 554 1042
rect 702 1038 706 1042
rect 846 1038 850 1042
rect 1406 1038 1410 1042
rect 1446 1038 1450 1042
rect 214 1028 218 1032
rect 1062 1027 1066 1031
rect 86 1018 90 1022
rect 126 1018 130 1022
rect 142 1018 146 1022
rect 182 1018 186 1022
rect 870 1018 874 1022
rect 1190 1018 1194 1022
rect 1254 1018 1258 1022
rect 482 1003 486 1007
rect 489 1003 493 1007
rect 22 988 26 992
rect 70 988 74 992
rect 166 988 170 992
rect 222 988 226 992
rect 294 988 298 992
rect 326 988 330 992
rect 462 988 466 992
rect 510 988 514 992
rect 566 988 570 992
rect 590 988 594 992
rect 622 988 626 992
rect 654 988 658 992
rect 694 988 698 992
rect 830 988 834 992
rect 854 988 858 992
rect 910 988 914 992
rect 1062 988 1066 992
rect 1158 988 1162 992
rect 1206 988 1210 992
rect 1254 988 1258 992
rect 1446 988 1450 992
rect 542 978 546 982
rect 14 968 18 972
rect 62 968 66 972
rect 158 968 162 972
rect 286 968 290 972
rect 318 968 322 972
rect 382 968 386 972
rect 390 968 394 972
rect 406 968 410 972
rect 438 968 442 972
rect 470 968 474 972
rect 518 968 522 972
rect 550 968 554 972
rect 598 968 602 972
rect 702 968 706 972
rect 782 968 786 972
rect 958 968 962 972
rect 966 968 970 972
rect 1430 968 1434 972
rect 1478 968 1482 972
rect 30 958 34 962
rect 78 958 82 962
rect 86 958 90 962
rect 14 948 18 952
rect 70 948 74 952
rect 174 958 178 962
rect 238 958 242 962
rect 302 958 306 962
rect 334 958 338 962
rect 374 958 378 962
rect 422 958 426 962
rect 454 958 458 962
rect 502 958 506 962
rect 534 958 538 962
rect 614 958 618 962
rect 686 958 690 962
rect 814 958 818 962
rect 894 958 898 962
rect 974 958 978 962
rect 990 958 994 962
rect 1022 958 1026 962
rect 1054 958 1058 962
rect 110 948 114 952
rect 142 948 146 952
rect 166 948 170 952
rect 182 948 186 952
rect 222 948 226 952
rect 270 948 274 952
rect 294 948 298 952
rect 326 948 330 952
rect 366 948 370 952
rect 382 948 386 952
rect 430 948 434 952
rect 462 948 466 952
rect 510 948 514 952
rect 542 948 546 952
rect 566 948 570 952
rect 606 948 610 952
rect 646 948 650 952
rect 678 948 682 952
rect 694 948 698 952
rect 742 948 746 952
rect 750 948 754 952
rect 766 948 770 952
rect 798 948 802 952
rect 830 948 834 952
rect 870 948 874 952
rect 910 948 914 952
rect 926 948 930 952
rect 966 948 970 952
rect 990 948 994 952
rect 1038 948 1042 952
rect 1054 948 1058 952
rect 1078 948 1082 952
rect 1102 948 1106 952
rect 1174 958 1178 962
rect 1254 958 1258 962
rect 1158 948 1162 952
rect 1182 948 1186 952
rect 1230 948 1234 952
rect 1270 948 1274 952
rect 1399 948 1403 952
rect 1406 948 1410 952
rect 1454 948 1458 952
rect 1462 948 1466 952
rect 38 938 42 942
rect 86 938 90 942
rect 118 938 122 942
rect 126 938 130 942
rect 134 938 138 942
rect 190 938 194 942
rect 262 938 266 942
rect 350 938 354 942
rect 358 938 362 942
rect 414 938 418 942
rect 638 938 642 942
rect 678 938 682 942
rect 718 938 722 942
rect 734 938 738 942
rect 750 938 754 942
rect 774 938 778 942
rect 806 938 810 942
rect 838 938 842 942
rect 886 938 890 942
rect 918 938 922 942
rect 982 938 986 942
rect 1030 938 1034 942
rect 1142 938 1146 942
rect 1190 938 1194 942
rect 1302 938 1306 942
rect 206 928 210 932
rect 246 928 250 932
rect 342 928 346 932
rect 582 928 586 932
rect 622 928 626 932
rect 654 928 658 932
rect 718 928 722 932
rect 926 928 930 932
rect 942 928 946 932
rect 1094 928 1098 932
rect 1118 928 1122 932
rect 1214 928 1218 932
rect 1318 928 1322 932
rect 1438 928 1442 932
rect 1486 928 1490 932
rect 46 918 50 922
rect 254 918 258 922
rect 1494 918 1498 922
rect 1002 903 1006 907
rect 1009 903 1013 907
rect 38 888 42 892
rect 78 888 82 892
rect 142 888 146 892
rect 222 888 226 892
rect 254 888 258 892
rect 438 888 442 892
rect 510 888 514 892
rect 590 888 594 892
rect 638 888 642 892
rect 670 888 674 892
rect 734 888 738 892
rect 790 888 794 892
rect 838 888 842 892
rect 846 888 850 892
rect 926 888 930 892
rect 1022 888 1026 892
rect 1062 888 1066 892
rect 1126 888 1130 892
rect 1246 888 1250 892
rect 1398 888 1402 892
rect 1414 888 1418 892
rect 30 878 34 882
rect 102 878 106 882
rect 374 878 378 882
rect 582 878 586 882
rect 870 878 874 882
rect 918 878 922 882
rect 950 878 954 882
rect 1174 878 1178 882
rect 1190 878 1194 882
rect 1198 878 1202 882
rect 1254 878 1258 882
rect 1406 878 1410 882
rect 1454 878 1458 882
rect 14 868 18 872
rect 62 868 66 872
rect 118 868 122 872
rect 182 868 186 872
rect 198 868 202 872
rect 246 868 250 872
rect 302 868 306 872
rect 334 868 338 872
rect 374 868 378 872
rect 390 868 394 872
rect 406 868 410 872
rect 422 868 426 872
rect 446 868 450 872
rect 478 868 482 872
rect 502 868 506 872
rect 526 868 530 872
rect 566 868 570 872
rect 574 868 578 872
rect 606 868 610 872
rect 614 868 618 872
rect 630 868 634 872
rect 662 868 666 872
rect 702 868 706 872
rect 718 868 722 872
rect 750 868 754 872
rect 758 868 762 872
rect 806 868 810 872
rect 854 868 858 872
rect 862 868 866 872
rect 886 868 890 872
rect 918 868 922 872
rect 934 868 938 872
rect 1054 868 1058 872
rect 1078 868 1082 872
rect 1102 868 1106 872
rect 1118 868 1122 872
rect 1166 868 1170 872
rect 1206 868 1210 872
rect 1230 868 1234 872
rect 1238 868 1242 872
rect 1262 868 1266 872
rect 1278 868 1282 872
rect 1294 868 1298 872
rect 1310 868 1314 872
rect 1326 868 1330 872
rect 1374 868 1378 872
rect 1390 868 1394 872
rect 1502 868 1506 872
rect 6 858 10 862
rect 54 858 58 862
rect 86 858 90 862
rect 102 858 106 862
rect 126 858 130 862
rect 150 858 154 862
rect 174 858 178 862
rect 254 858 258 862
rect 270 858 274 862
rect 286 858 290 862
rect 302 858 306 862
rect 326 858 330 862
rect 358 858 362 862
rect 398 858 402 862
rect 446 858 450 862
rect 478 858 482 862
rect 526 858 530 862
rect 558 858 562 862
rect 654 858 658 862
rect 694 858 698 862
rect 822 858 826 862
rect 894 858 898 862
rect 966 858 970 862
rect 1110 858 1114 862
rect 1166 858 1170 862
rect 1230 858 1234 862
rect 1270 858 1274 862
rect 1286 858 1290 862
rect 1302 858 1306 862
rect 1358 858 1362 862
rect 1382 858 1386 862
rect 1430 858 1434 862
rect 1462 858 1466 862
rect 38 848 42 852
rect 94 848 98 852
rect 158 848 162 852
rect 166 848 170 852
rect 278 848 282 852
rect 310 848 314 852
rect 342 848 346 852
rect 366 848 370 852
rect 406 848 410 852
rect 430 848 434 852
rect 454 848 458 852
rect 518 848 522 852
rect 550 848 554 852
rect 590 848 594 852
rect 614 848 618 852
rect 638 848 642 852
rect 670 848 674 852
rect 726 848 730 852
rect 734 848 738 852
rect 910 848 914 852
rect 1062 848 1066 852
rect 1142 848 1146 852
rect 1286 848 1290 852
rect 1318 848 1322 852
rect 1414 848 1418 852
rect 1486 848 1490 852
rect 78 838 82 842
rect 158 838 162 842
rect 182 838 186 842
rect 326 838 330 842
rect 350 838 354 842
rect 534 838 538 842
rect 1478 838 1482 842
rect 30 818 34 822
rect 846 818 850 822
rect 1094 818 1098 822
rect 1494 818 1498 822
rect 482 803 486 807
rect 489 803 493 807
rect 22 788 26 792
rect 158 788 162 792
rect 502 788 506 792
rect 550 788 554 792
rect 606 788 610 792
rect 646 788 650 792
rect 670 788 674 792
rect 702 788 706 792
rect 726 788 730 792
rect 774 788 778 792
rect 822 788 826 792
rect 878 788 882 792
rect 1038 788 1042 792
rect 1110 788 1114 792
rect 1190 788 1194 792
rect 1414 788 1418 792
rect 1462 788 1466 792
rect 430 778 434 782
rect 526 778 530 782
rect 582 778 586 782
rect 1286 778 1290 782
rect 14 768 18 772
rect 78 768 82 772
rect 150 768 154 772
rect 422 768 426 772
rect 510 768 514 772
rect 558 768 562 772
rect 590 768 594 772
rect 766 768 770 772
rect 1374 768 1378 772
rect 30 758 34 762
rect 70 758 74 762
rect 94 758 98 762
rect 134 758 138 762
rect 166 758 170 762
rect 198 758 202 762
rect 214 758 218 762
rect 246 758 250 762
rect 22 748 26 752
rect 38 748 42 752
rect 54 748 58 752
rect 86 748 90 752
rect 102 748 106 752
rect 126 748 130 752
rect 142 748 146 752
rect 198 748 202 752
rect 230 748 234 752
rect 278 758 282 762
rect 334 758 338 762
rect 350 758 354 762
rect 358 758 362 762
rect 438 758 442 762
rect 494 758 498 762
rect 534 758 538 762
rect 574 758 578 762
rect 630 758 634 762
rect 686 758 690 762
rect 742 758 746 762
rect 782 758 786 762
rect 830 758 834 762
rect 862 758 866 762
rect 918 758 922 762
rect 942 758 946 762
rect 294 748 298 752
rect 334 748 338 752
rect 406 748 410 752
rect 430 748 434 752
rect 470 748 474 752
rect 502 748 506 752
rect 550 748 554 752
rect 582 748 586 752
rect 606 748 610 752
rect 646 748 650 752
rect 710 748 714 752
rect 726 748 730 752
rect 862 748 866 752
rect 902 748 906 752
rect 958 748 962 752
rect 1014 748 1018 752
rect 1078 748 1082 752
rect 1086 748 1090 752
rect 1134 748 1138 752
rect 1150 748 1154 752
rect 1190 748 1194 752
rect 1198 748 1202 752
rect 1214 758 1218 762
rect 1326 758 1330 762
rect 1358 758 1362 762
rect 1390 758 1394 762
rect 1398 758 1402 762
rect 1502 758 1506 762
rect 1254 748 1258 752
rect 1270 748 1274 752
rect 1294 748 1298 752
rect 1342 748 1346 752
rect 1358 748 1362 752
rect 1374 748 1378 752
rect 1414 748 1418 752
rect 1454 748 1458 752
rect 46 738 50 742
rect 62 738 66 742
rect 118 738 122 742
rect 182 738 186 742
rect 190 738 194 742
rect 222 738 226 742
rect 270 738 274 742
rect 318 738 322 742
rect 374 738 378 742
rect 382 738 386 742
rect 398 738 402 742
rect 462 738 466 742
rect 662 738 666 742
rect 718 738 722 742
rect 750 738 754 742
rect 766 738 770 742
rect 790 738 794 742
rect 806 738 810 742
rect 814 738 818 742
rect 830 738 834 742
rect 838 738 842 742
rect 870 738 874 742
rect 894 738 898 742
rect 926 738 930 742
rect 942 738 946 742
rect 950 738 954 742
rect 990 738 994 742
rect 1030 738 1034 742
rect 1070 738 1074 742
rect 1086 738 1090 742
rect 1142 738 1146 742
rect 1222 738 1226 742
rect 1246 738 1250 742
rect 1262 738 1266 742
rect 1294 738 1298 742
rect 1318 738 1322 742
rect 1334 738 1338 742
rect 1366 738 1370 742
rect 1422 738 1426 742
rect 1438 738 1442 742
rect 1470 738 1474 742
rect 102 728 106 732
rect 174 728 178 732
rect 262 728 266 732
rect 278 728 282 732
rect 382 728 386 732
rect 446 728 450 732
rect 454 728 458 732
rect 534 728 538 732
rect 622 728 626 732
rect 694 728 698 732
rect 886 728 890 732
rect 1046 728 1050 732
rect 1054 728 1058 732
rect 1110 728 1114 732
rect 1166 728 1170 732
rect 1230 728 1234 732
rect 1430 728 1434 732
rect 358 718 362 722
rect 782 718 786 722
rect 798 718 802 722
rect 918 718 922 722
rect 990 718 994 722
rect 1062 718 1066 722
rect 1102 718 1106 722
rect 1118 718 1122 722
rect 1238 718 1242 722
rect 1462 718 1466 722
rect 1486 718 1490 722
rect 1002 703 1006 707
rect 1009 703 1013 707
rect 46 688 50 692
rect 110 688 114 692
rect 126 688 130 692
rect 166 688 170 692
rect 230 688 234 692
rect 318 688 322 692
rect 342 688 346 692
rect 366 688 370 692
rect 390 688 394 692
rect 446 688 450 692
rect 454 688 458 692
rect 526 688 530 692
rect 534 688 538 692
rect 646 688 650 692
rect 686 688 690 692
rect 710 688 714 692
rect 734 688 738 692
rect 846 688 850 692
rect 870 688 874 692
rect 958 688 962 692
rect 1054 688 1058 692
rect 1142 688 1146 692
rect 1302 688 1306 692
rect 1430 688 1434 692
rect 1438 688 1442 692
rect 30 678 34 682
rect 14 668 18 672
rect 54 678 58 682
rect 238 678 242 682
rect 310 678 314 682
rect 606 678 610 682
rect 638 678 642 682
rect 694 678 698 682
rect 878 678 882 682
rect 902 678 906 682
rect 950 678 954 682
rect 982 678 986 682
rect 990 678 994 682
rect 1150 678 1154 682
rect 1190 678 1194 682
rect 1222 678 1226 682
rect 1270 678 1274 682
rect 1310 678 1314 682
rect 1318 678 1322 682
rect 78 668 82 672
rect 214 668 218 672
rect 238 668 242 672
rect 278 668 282 672
rect 286 668 290 672
rect 302 668 306 672
rect 326 668 330 672
rect 366 668 370 672
rect 382 668 386 672
rect 422 668 426 672
rect 502 668 506 672
rect 550 668 554 672
rect 558 668 562 672
rect 574 668 578 672
rect 598 668 602 672
rect 606 668 610 672
rect 622 668 626 672
rect 654 668 658 672
rect 678 668 682 672
rect 702 668 706 672
rect 742 668 746 672
rect 750 668 754 672
rect 822 668 826 672
rect 854 668 858 672
rect 1014 668 1018 672
rect 1046 668 1050 672
rect 1094 668 1098 672
rect 1126 668 1130 672
rect 1150 668 1154 672
rect 1174 668 1178 672
rect 1214 668 1218 672
rect 1238 668 1242 672
rect 1262 668 1266 672
rect 1286 668 1290 672
rect 1334 668 1338 672
rect 1350 668 1354 672
rect 1374 668 1378 672
rect 1390 668 1394 672
rect 1454 668 1458 672
rect 1470 678 1474 682
rect 1486 668 1490 672
rect 6 658 10 662
rect 86 658 90 662
rect 102 658 106 662
rect 142 658 146 662
rect 166 658 170 662
rect 190 658 194 662
rect 206 658 210 662
rect 222 658 226 662
rect 254 658 258 662
rect 270 658 274 662
rect 334 658 338 662
rect 430 658 434 662
rect 510 658 514 662
rect 566 658 570 662
rect 582 658 586 662
rect 598 658 602 662
rect 630 658 634 662
rect 662 658 666 662
rect 670 658 674 662
rect 750 658 754 662
rect 774 658 778 662
rect 790 658 794 662
rect 814 658 818 662
rect 894 658 898 662
rect 918 658 922 662
rect 926 658 930 662
rect 966 658 970 662
rect 974 658 978 662
rect 1022 658 1026 662
rect 1046 658 1050 662
rect 1118 658 1122 662
rect 1126 658 1130 662
rect 1166 658 1170 662
rect 1206 658 1210 662
rect 1254 658 1258 662
rect 1270 658 1274 662
rect 1326 658 1330 662
rect 1342 658 1346 662
rect 1358 658 1362 662
rect 1366 658 1370 662
rect 1398 658 1402 662
rect 1414 658 1418 662
rect 1494 658 1498 662
rect 94 648 98 652
rect 150 648 154 652
rect 158 648 162 652
rect 286 648 290 652
rect 342 648 346 652
rect 366 648 370 652
rect 390 648 394 652
rect 454 648 458 652
rect 526 648 530 652
rect 534 648 538 652
rect 718 648 722 652
rect 774 648 778 652
rect 846 648 850 652
rect 870 648 874 652
rect 902 648 906 652
rect 942 648 946 652
rect 1038 648 1042 652
rect 1062 648 1066 652
rect 1070 648 1074 652
rect 1102 648 1106 652
rect 1182 648 1186 652
rect 1230 648 1234 652
rect 1238 648 1242 652
rect 1302 648 1306 652
rect 1374 648 1378 652
rect 1406 648 1410 652
rect 110 638 114 642
rect 166 638 170 642
rect 1422 638 1426 642
rect 254 628 258 632
rect 758 618 762 622
rect 806 618 810 622
rect 926 618 930 622
rect 1086 618 1090 622
rect 482 603 486 607
rect 489 603 493 607
rect 134 588 138 592
rect 190 588 194 592
rect 214 588 218 592
rect 350 588 354 592
rect 494 588 498 592
rect 558 588 562 592
rect 574 588 578 592
rect 614 588 618 592
rect 638 588 642 592
rect 1166 588 1170 592
rect 1358 588 1362 592
rect 1446 588 1450 592
rect 246 578 250 582
rect 318 578 322 582
rect 38 568 42 572
rect 54 568 58 572
rect 86 568 90 572
rect 118 568 122 572
rect 198 568 202 572
rect 222 568 226 572
rect 254 568 258 572
rect 326 568 330 572
rect 358 568 362 572
rect 790 568 794 572
rect 822 568 826 572
rect 1302 568 1306 572
rect 1350 568 1354 572
rect 30 548 34 552
rect 182 558 186 562
rect 238 558 242 562
rect 270 558 274 562
rect 310 558 314 562
rect 342 558 346 562
rect 622 558 626 562
rect 774 558 778 562
rect 806 558 810 562
rect 878 558 882 562
rect 926 558 930 562
rect 958 558 962 562
rect 1014 558 1018 562
rect 1134 558 1138 562
rect 1182 558 1186 562
rect 1206 558 1210 562
rect 1222 558 1226 562
rect 1294 558 1298 562
rect 1334 558 1338 562
rect 134 548 138 552
rect 150 548 154 552
rect 190 548 194 552
rect 230 548 234 552
rect 262 548 266 552
rect 302 548 306 552
rect 318 548 322 552
rect 350 548 354 552
rect 382 548 386 552
rect 398 548 402 552
rect 414 548 418 552
rect 430 548 434 552
rect 446 548 450 552
rect 510 548 514 552
rect 542 548 546 552
rect 566 548 570 552
rect 598 548 602 552
rect 686 548 690 552
rect 734 548 738 552
rect 790 548 794 552
rect 830 548 834 552
rect 862 548 866 552
rect 886 548 890 552
rect 910 548 914 552
rect 942 548 946 552
rect 966 548 970 552
rect 982 548 986 552
rect 1014 548 1018 552
rect 1054 548 1058 552
rect 1070 548 1074 552
rect 1102 548 1106 552
rect 1118 548 1122 552
rect 1166 548 1170 552
rect 1214 548 1218 552
rect 1238 548 1242 552
rect 1278 548 1282 552
rect 1326 548 1330 552
rect 1342 548 1346 552
rect 1390 548 1394 552
rect 1446 548 1450 552
rect 1462 548 1466 552
rect 1502 548 1506 552
rect 70 538 74 542
rect 110 538 114 542
rect 142 538 146 542
rect 158 538 162 542
rect 294 538 298 542
rect 374 538 378 542
rect 390 538 394 542
rect 414 538 418 542
rect 422 538 426 542
rect 438 538 442 542
rect 470 538 474 542
rect 510 538 514 542
rect 534 538 538 542
rect 590 538 594 542
rect 606 538 610 542
rect 630 538 634 542
rect 766 538 770 542
rect 798 538 802 542
rect 854 538 858 542
rect 902 538 906 542
rect 934 538 938 542
rect 1006 538 1010 542
rect 1054 538 1058 542
rect 1094 538 1098 542
rect 1110 538 1114 542
rect 1158 538 1162 542
rect 1190 538 1194 542
rect 1246 538 1250 542
rect 1270 538 1274 542
rect 1318 538 1322 542
rect 1366 538 1370 542
rect 1382 538 1386 542
rect 1414 538 1418 542
rect 1422 538 1426 542
rect 6 528 10 532
rect 78 528 82 532
rect 174 528 178 532
rect 278 528 282 532
rect 422 528 426 532
rect 454 528 458 532
rect 462 528 466 532
rect 518 528 522 532
rect 550 528 554 532
rect 574 528 578 532
rect 670 528 674 532
rect 694 528 698 532
rect 710 528 714 532
rect 750 528 754 532
rect 846 528 850 532
rect 1038 528 1042 532
rect 1054 528 1058 532
rect 1078 528 1082 532
rect 1230 528 1234 532
rect 1254 528 1258 532
rect 1262 528 1266 532
rect 1422 528 1426 532
rect 1462 528 1466 532
rect 1478 528 1482 532
rect 1486 528 1490 532
rect 38 518 42 522
rect 86 518 90 522
rect 166 518 170 522
rect 286 518 290 522
rect 638 518 642 522
rect 678 518 682 522
rect 758 518 762 522
rect 838 518 842 522
rect 894 518 898 522
rect 926 518 930 522
rect 1086 518 1090 522
rect 1150 518 1154 522
rect 1198 518 1202 522
rect 1374 518 1378 522
rect 1494 518 1498 522
rect 1002 503 1006 507
rect 1009 503 1013 507
rect 62 488 66 492
rect 102 488 106 492
rect 254 488 258 492
rect 374 488 378 492
rect 534 488 538 492
rect 574 488 578 492
rect 614 488 618 492
rect 646 488 650 492
rect 702 488 706 492
rect 1046 488 1050 492
rect 1134 488 1138 492
rect 1382 488 1386 492
rect 1414 488 1418 492
rect 1494 488 1498 492
rect 166 478 170 482
rect 182 478 186 482
rect 246 478 250 482
rect 422 478 426 482
rect 430 478 434 482
rect 502 478 506 482
rect 798 478 802 482
rect 1118 478 1122 482
rect 1126 478 1130 482
rect 1262 478 1266 482
rect 1350 478 1354 482
rect 1486 478 1490 482
rect 22 466 26 470
rect 30 468 34 472
rect 38 468 42 472
rect 54 468 58 472
rect 94 468 98 472
rect 190 468 194 472
rect 238 468 242 472
rect 262 468 266 472
rect 302 468 306 472
rect 318 468 322 472
rect 342 468 346 472
rect 358 468 362 472
rect 398 468 402 472
rect 430 468 434 472
rect 446 468 450 472
rect 462 468 466 472
rect 478 468 482 472
rect 494 468 498 472
rect 518 468 522 472
rect 550 468 554 472
rect 558 468 562 472
rect 574 468 578 472
rect 606 468 610 472
rect 702 468 706 472
rect 718 468 722 472
rect 726 468 730 472
rect 742 468 746 472
rect 774 468 778 472
rect 806 468 810 472
rect 822 468 826 472
rect 838 468 842 472
rect 878 468 882 472
rect 894 468 898 472
rect 902 468 906 472
rect 934 468 938 472
rect 78 458 82 462
rect 142 458 146 462
rect 166 458 170 462
rect 270 458 274 462
rect 294 458 298 462
rect 350 458 354 462
rect 390 458 394 462
rect 406 458 410 462
rect 454 458 458 462
rect 526 458 530 462
rect 598 458 602 462
rect 662 458 666 462
rect 766 458 770 462
rect 782 458 786 462
rect 790 458 794 462
rect 814 458 818 462
rect 830 458 834 462
rect 846 458 850 462
rect 854 458 858 462
rect 886 458 890 462
rect 910 458 914 462
rect 958 468 962 472
rect 1006 468 1010 472
rect 1038 468 1042 472
rect 1070 468 1074 472
rect 1078 468 1082 472
rect 1182 468 1186 472
rect 1206 468 1210 472
rect 1230 468 1234 472
rect 1246 468 1250 472
rect 1262 468 1266 472
rect 1294 468 1298 472
rect 1342 468 1346 472
rect 1398 468 1402 472
rect 1406 468 1410 472
rect 1478 468 1482 472
rect 998 458 1002 462
rect 1014 458 1018 462
rect 1030 458 1034 462
rect 1062 458 1066 462
rect 1086 458 1090 462
rect 1150 458 1154 462
rect 1158 458 1162 462
rect 1190 458 1194 462
rect 1214 458 1218 462
rect 1238 458 1242 462
rect 1270 458 1274 462
rect 1286 458 1290 462
rect 1310 458 1314 462
rect 1366 458 1370 462
rect 1398 458 1402 462
rect 1502 458 1506 462
rect 54 448 58 452
rect 86 448 90 452
rect 110 448 114 452
rect 142 448 146 452
rect 158 448 162 452
rect 278 448 282 452
rect 310 448 314 452
rect 366 448 370 452
rect 462 448 466 452
rect 534 448 538 452
rect 574 448 578 452
rect 582 448 586 452
rect 614 448 618 452
rect 702 448 706 452
rect 726 448 730 452
rect 742 448 746 452
rect 830 448 834 452
rect 862 448 866 452
rect 870 448 874 452
rect 934 448 938 452
rect 950 448 954 452
rect 990 448 994 452
rect 1046 448 1050 452
rect 1102 448 1106 452
rect 1174 448 1178 452
rect 1206 448 1210 452
rect 1214 448 1218 452
rect 1270 448 1274 452
rect 1302 448 1306 452
rect 1318 448 1322 452
rect 1430 448 1434 452
rect 1454 448 1458 452
rect 78 438 82 442
rect 406 438 410 442
rect 1366 438 1370 442
rect 6 418 10 422
rect 214 418 218 422
rect 622 418 626 422
rect 686 418 690 422
rect 710 418 714 422
rect 734 418 738 422
rect 766 418 770 422
rect 1022 418 1026 422
rect 1086 418 1090 422
rect 1110 418 1114 422
rect 1158 418 1162 422
rect 1310 418 1314 422
rect 1334 418 1338 422
rect 482 403 486 407
rect 489 403 493 407
rect 22 388 26 392
rect 78 388 82 392
rect 110 388 114 392
rect 142 388 146 392
rect 206 388 210 392
rect 310 388 314 392
rect 342 388 346 392
rect 366 388 370 392
rect 398 388 402 392
rect 614 388 618 392
rect 742 388 746 392
rect 758 388 762 392
rect 854 388 858 392
rect 1286 388 1290 392
rect 1334 388 1338 392
rect 1366 388 1370 392
rect 1414 388 1418 392
rect 574 378 578 382
rect 1054 378 1058 382
rect 1086 378 1090 382
rect 86 368 90 372
rect 150 368 154 372
rect 214 368 218 372
rect 422 368 426 372
rect 774 368 778 372
rect 886 368 890 372
rect 1046 368 1050 372
rect 1358 368 1362 372
rect 6 358 10 362
rect 70 358 74 362
rect 126 358 130 362
rect 134 358 138 362
rect 198 358 202 362
rect 246 358 250 362
rect 286 358 290 362
rect 358 358 362 362
rect 454 358 458 362
rect 710 358 714 362
rect 22 348 26 352
rect 38 348 42 352
rect 78 348 82 352
rect 110 348 114 352
rect 142 348 146 352
rect 846 358 850 362
rect 974 358 978 362
rect 1030 358 1034 362
rect 1070 358 1074 362
rect 1182 358 1186 362
rect 1206 358 1210 362
rect 1374 358 1378 362
rect 1438 358 1442 362
rect 206 348 210 352
rect 326 348 330 352
rect 382 348 386 352
rect 30 338 34 342
rect 46 338 50 342
rect 54 338 58 342
rect 102 338 106 342
rect 166 338 170 342
rect 182 338 186 342
rect 230 338 234 342
rect 278 338 282 342
rect 302 338 306 342
rect 374 338 378 342
rect 446 348 450 352
rect 526 348 530 352
rect 558 348 562 352
rect 590 348 594 352
rect 598 348 602 352
rect 646 348 650 352
rect 670 348 674 352
rect 686 348 690 352
rect 694 348 698 352
rect 702 348 706 352
rect 718 348 722 352
rect 758 348 762 352
rect 798 348 802 352
rect 822 348 826 352
rect 838 348 842 352
rect 886 348 890 352
rect 902 348 906 352
rect 918 348 922 352
rect 926 348 930 352
rect 958 348 962 352
rect 1014 348 1018 352
rect 1094 348 1098 352
rect 1102 348 1106 352
rect 1134 348 1138 352
rect 1158 348 1162 352
rect 1190 348 1194 352
rect 1246 348 1250 352
rect 1366 348 1370 352
rect 1382 348 1386 352
rect 1414 348 1418 352
rect 1438 348 1442 352
rect 422 338 426 342
rect 438 338 442 342
rect 454 338 458 342
rect 470 338 474 342
rect 478 338 482 342
rect 550 338 554 342
rect 686 338 690 342
rect 718 338 722 342
rect 750 338 754 342
rect 806 338 810 342
rect 814 338 818 342
rect 862 338 866 342
rect 910 338 914 342
rect 1022 338 1026 342
rect 1046 338 1050 342
rect 1062 338 1066 342
rect 1094 338 1098 342
rect 1118 338 1122 342
rect 1126 338 1130 342
rect 1158 338 1162 342
rect 1190 338 1194 342
rect 1222 338 1226 342
rect 1318 338 1322 342
rect 1342 338 1346 342
rect 1398 338 1402 342
rect 1454 338 1458 342
rect 1486 338 1490 342
rect 62 328 66 332
rect 166 328 170 332
rect 318 328 322 332
rect 366 328 370 332
rect 662 328 666 332
rect 742 328 746 332
rect 838 328 842 332
rect 870 328 874 332
rect 894 328 898 332
rect 942 328 946 332
rect 982 328 986 332
rect 1118 328 1122 332
rect 1214 328 1218 332
rect 1270 328 1274 332
rect 1326 328 1330 332
rect 1414 328 1418 332
rect 1430 328 1434 332
rect 1486 328 1490 332
rect 286 318 290 322
rect 454 318 458 322
rect 782 318 786 322
rect 974 318 978 322
rect 990 318 994 322
rect 1150 318 1154 322
rect 1182 318 1186 322
rect 1462 318 1466 322
rect 1002 303 1006 307
rect 1009 303 1013 307
rect 70 288 74 292
rect 110 288 114 292
rect 150 288 154 292
rect 190 288 194 292
rect 518 288 522 292
rect 630 288 634 292
rect 710 288 714 292
rect 742 288 746 292
rect 798 288 802 292
rect 822 288 826 292
rect 862 288 866 292
rect 958 288 962 292
rect 1038 288 1042 292
rect 1110 288 1114 292
rect 1174 288 1178 292
rect 1382 288 1386 292
rect 1406 288 1410 292
rect 1502 288 1506 292
rect 118 278 122 282
rect 622 278 626 282
rect 646 278 650 282
rect 782 278 786 282
rect 790 278 794 282
rect 830 278 834 282
rect 934 278 938 282
rect 966 278 970 282
rect 1054 278 1058 282
rect 1118 278 1122 282
rect 1142 278 1146 282
rect 1150 278 1154 282
rect 1182 278 1186 282
rect 1326 278 1330 282
rect 1390 278 1394 282
rect 1438 278 1442 282
rect 1454 278 1458 282
rect 1478 278 1482 282
rect 1486 278 1490 282
rect 6 268 10 272
rect 54 268 58 272
rect 102 268 106 272
rect 142 268 146 272
rect 158 268 162 272
rect 206 268 210 272
rect 222 268 226 272
rect 294 268 298 272
rect 350 268 354 272
rect 390 268 394 272
rect 462 268 466 272
rect 526 268 530 272
rect 534 268 538 272
rect 582 268 586 272
rect 654 268 658 272
rect 686 268 690 272
rect 694 268 698 272
rect 814 268 818 272
rect 838 268 842 272
rect 878 268 882 272
rect 950 268 954 272
rect 974 268 978 272
rect 998 268 1002 272
rect 1014 268 1018 272
rect 1022 266 1026 270
rect 1086 268 1090 272
rect 1102 268 1106 272
rect 1134 268 1138 272
rect 1166 268 1170 272
rect 1182 268 1186 272
rect 1214 268 1218 272
rect 1246 268 1250 272
rect 1286 268 1290 272
rect 1302 268 1306 272
rect 1334 268 1338 272
rect 1374 268 1378 272
rect 1414 268 1418 272
rect 1430 268 1434 272
rect 78 258 82 262
rect 94 258 98 262
rect 166 258 170 262
rect 182 258 186 262
rect 222 258 226 262
rect 246 258 250 262
rect 278 258 282 262
rect 326 258 330 262
rect 366 258 370 262
rect 382 258 386 262
rect 414 258 418 262
rect 438 258 442 262
rect 502 258 506 262
rect 566 258 570 262
rect 582 258 586 262
rect 606 258 610 262
rect 662 258 666 262
rect 678 258 682 262
rect 710 258 714 262
rect 750 258 754 262
rect 758 258 762 262
rect 766 258 770 262
rect 806 258 810 262
rect 846 258 850 262
rect 894 258 898 262
rect 918 258 922 262
rect 926 258 930 262
rect 942 258 946 262
rect 1078 258 1082 262
rect 1094 258 1098 262
rect 1126 258 1130 262
rect 1158 258 1162 262
rect 1238 258 1242 262
rect 1262 258 1266 262
rect 1278 258 1282 262
rect 1310 258 1314 262
rect 1326 258 1330 262
rect 1414 258 1418 262
rect 1462 258 1466 262
rect 86 248 90 252
rect 174 248 178 252
rect 254 248 258 252
rect 286 248 290 252
rect 342 248 346 252
rect 422 248 426 252
rect 430 248 434 252
rect 550 248 554 252
rect 590 248 594 252
rect 638 248 642 252
rect 654 248 658 252
rect 710 248 714 252
rect 862 248 866 252
rect 870 248 874 252
rect 990 248 994 252
rect 1054 248 1058 252
rect 1078 248 1082 252
rect 1190 248 1194 252
rect 1222 248 1226 252
rect 1358 248 1362 252
rect 38 238 42 242
rect 86 238 90 242
rect 190 238 194 242
rect 238 238 242 242
rect 270 238 274 242
rect 406 238 410 242
rect 446 238 450 242
rect 246 218 250 222
rect 278 218 282 222
rect 366 218 370 222
rect 398 218 402 222
rect 438 218 442 222
rect 774 218 778 222
rect 1046 218 1050 222
rect 482 203 486 207
rect 489 203 493 207
rect 22 188 26 192
rect 86 188 90 192
rect 198 188 202 192
rect 598 188 602 192
rect 798 188 802 192
rect 934 188 938 192
rect 1230 188 1234 192
rect 1262 188 1266 192
rect 1462 188 1466 192
rect 150 178 154 182
rect 14 168 18 172
rect 46 168 50 172
rect 206 168 210 172
rect 742 178 746 182
rect 246 168 250 172
rect 342 168 346 172
rect 358 168 362 172
rect 742 168 746 172
rect 1054 168 1058 172
rect 1070 168 1074 172
rect 1158 168 1162 172
rect 1198 168 1202 172
rect 1278 168 1282 172
rect 1334 168 1338 172
rect 30 158 34 162
rect 62 158 66 162
rect 70 158 74 162
rect 134 158 138 162
rect 190 158 194 162
rect 230 158 234 162
rect 310 158 314 162
rect 374 158 378 162
rect 558 158 562 162
rect 726 158 730 162
rect 766 158 770 162
rect 862 158 866 162
rect 942 158 946 162
rect 1310 158 1314 162
rect 1318 158 1322 162
rect 1382 158 1386 162
rect 22 148 26 152
rect 38 148 42 152
rect 54 148 58 152
rect 126 148 130 152
rect 174 148 178 152
rect 182 148 186 152
rect 214 148 218 152
rect 238 148 242 152
rect 286 148 290 152
rect 326 148 330 152
rect 350 148 354 152
rect 366 148 370 152
rect 406 148 410 152
rect 430 148 434 152
rect 486 148 490 152
rect 510 148 514 152
rect 542 148 546 152
rect 582 148 586 152
rect 606 148 610 152
rect 614 148 618 152
rect 638 148 642 152
rect 670 148 674 152
rect 678 148 682 152
rect 694 148 698 152
rect 726 148 730 152
rect 734 148 738 152
rect 750 148 754 152
rect 798 148 802 152
rect 862 148 866 152
rect 878 148 882 152
rect 94 138 98 142
rect 118 138 122 142
rect 158 138 162 142
rect 278 138 282 142
rect 294 138 298 142
rect 318 138 322 142
rect 398 138 402 142
rect 414 138 418 142
rect 454 138 458 142
rect 478 138 482 142
rect 518 138 522 142
rect 662 138 666 142
rect 702 138 706 142
rect 958 148 962 152
rect 990 148 994 152
rect 1014 148 1018 152
rect 1046 148 1050 152
rect 1054 148 1058 152
rect 1070 148 1074 152
rect 1102 148 1106 152
rect 1118 148 1122 152
rect 1134 148 1138 152
rect 1150 148 1154 152
rect 1190 148 1194 152
rect 1206 148 1210 152
rect 1270 148 1274 152
rect 1286 148 1290 152
rect 1334 148 1338 152
rect 1350 148 1354 152
rect 1366 148 1370 152
rect 1382 148 1386 152
rect 1398 148 1402 152
rect 1438 148 1442 152
rect 1478 148 1482 152
rect 1486 148 1490 152
rect 854 138 858 142
rect 886 138 890 142
rect 894 138 898 142
rect 902 138 906 142
rect 910 138 914 142
rect 918 138 922 142
rect 998 138 1002 142
rect 1046 138 1050 142
rect 1078 138 1082 142
rect 1094 138 1098 142
rect 1110 138 1114 142
rect 1142 138 1146 142
rect 1206 138 1210 142
rect 1262 138 1266 142
rect 1286 138 1290 142
rect 1350 138 1354 142
rect 1374 138 1378 142
rect 1406 138 1410 142
rect 1422 138 1426 142
rect 102 128 106 132
rect 262 128 266 132
rect 382 128 386 132
rect 414 128 418 132
rect 462 128 466 132
rect 534 128 538 132
rect 622 128 626 132
rect 638 128 642 132
rect 654 128 658 132
rect 766 128 770 132
rect 782 128 786 132
rect 1022 128 1026 132
rect 1166 128 1170 132
rect 1246 128 1250 132
rect 1310 128 1314 132
rect 1350 128 1354 132
rect 1430 128 1434 132
rect 1502 128 1506 132
rect 270 118 274 122
rect 302 118 306 122
rect 390 118 394 122
rect 470 118 474 122
rect 526 118 530 122
rect 686 118 690 122
rect 862 118 866 122
rect 1118 118 1122 122
rect 1174 118 1178 122
rect 1002 103 1006 107
rect 1009 103 1013 107
rect 30 88 34 92
rect 78 88 82 92
rect 126 88 130 92
rect 206 88 210 92
rect 246 88 250 92
rect 254 88 258 92
rect 494 88 498 92
rect 582 88 586 92
rect 614 88 618 92
rect 646 88 650 92
rect 662 88 666 92
rect 718 88 722 92
rect 830 88 834 92
rect 870 88 874 92
rect 958 88 962 92
rect 1094 88 1098 92
rect 1190 88 1194 92
rect 1414 88 1418 92
rect 1446 88 1450 92
rect 166 78 170 82
rect 238 78 242 82
rect 350 78 354 82
rect 54 68 58 72
rect 62 68 66 72
rect 118 68 122 72
rect 174 68 178 72
rect 182 68 186 72
rect 230 68 234 72
rect 278 68 282 72
rect 286 68 290 72
rect 334 68 338 72
rect 358 68 362 72
rect 374 68 378 72
rect 446 68 450 72
rect 654 78 658 82
rect 694 78 698 82
rect 734 78 738 82
rect 782 78 786 82
rect 822 78 826 82
rect 846 78 850 82
rect 862 78 866 82
rect 1046 78 1050 82
rect 1110 78 1114 82
rect 1150 78 1154 82
rect 1166 78 1170 82
rect 1230 78 1234 82
rect 1278 78 1282 82
rect 1342 78 1346 82
rect 1366 78 1370 82
rect 1422 78 1426 82
rect 1454 78 1458 82
rect 470 68 474 72
rect 534 68 538 72
rect 566 68 570 72
rect 574 68 578 72
rect 678 68 682 72
rect 726 68 730 72
rect 758 68 762 72
rect 790 68 794 72
rect 910 68 914 72
rect 926 68 930 72
rect 942 68 946 72
rect 950 68 954 72
rect 982 68 986 72
rect 1006 68 1010 72
rect 1022 68 1026 72
rect 1126 68 1130 72
rect 1158 68 1162 72
rect 1174 68 1178 72
rect 1222 68 1226 72
rect 1230 68 1234 72
rect 1246 68 1250 72
rect 1294 68 1298 72
rect 1326 68 1330 72
rect 1374 68 1378 72
rect 1438 68 1442 72
rect 1462 68 1466 72
rect 1478 68 1482 72
rect 150 58 154 62
rect 270 58 274 62
rect 366 58 370 62
rect 478 58 482 62
rect 494 58 498 62
rect 542 58 546 62
rect 598 58 602 62
rect 670 58 674 62
rect 702 58 706 62
rect 734 58 738 62
rect 750 58 754 62
rect 798 58 802 62
rect 846 58 850 62
rect 862 58 866 62
rect 886 58 890 62
rect 902 58 906 62
rect 934 58 938 62
rect 958 58 962 62
rect 990 58 994 62
rect 1014 58 1018 62
rect 1030 58 1034 62
rect 1062 58 1066 62
rect 1102 58 1106 62
rect 1118 58 1122 62
rect 1150 58 1154 62
rect 1198 58 1202 62
rect 1214 58 1218 62
rect 1254 58 1258 62
rect 1302 58 1306 62
rect 1326 58 1330 62
rect 1398 58 1402 62
rect 1430 58 1434 62
rect 1470 58 1474 62
rect 254 48 258 52
rect 302 48 306 52
rect 398 48 402 52
rect 646 48 650 52
rect 782 48 786 52
rect 798 48 802 52
rect 814 48 818 52
rect 1030 48 1034 52
rect 1078 48 1082 52
rect 1198 48 1202 52
rect 1270 48 1274 52
rect 1318 48 1322 52
rect 1494 48 1498 52
rect 518 38 522 42
rect 590 38 594 42
rect 482 3 486 7
rect 489 3 493 7
<< metal2 >>
rect 774 1328 778 1332
rect 910 1328 914 1332
rect 466 1288 470 1291
rect 42 1268 46 1271
rect 6 1262 9 1268
rect 14 1242 17 1268
rect 22 1242 25 1258
rect 14 1231 17 1238
rect 14 1228 25 1231
rect 22 1192 25 1228
rect 30 1212 33 1248
rect 38 1242 41 1258
rect 62 1212 65 1278
rect 70 1272 73 1278
rect 86 1252 89 1268
rect 94 1262 97 1268
rect 102 1252 105 1288
rect 774 1282 777 1328
rect 910 1282 913 1328
rect 1502 1318 1518 1321
rect 1000 1303 1002 1307
rect 1006 1303 1009 1307
rect 1013 1303 1016 1307
rect 570 1278 574 1281
rect 658 1278 662 1281
rect 1210 1278 1214 1281
rect 1378 1278 1382 1281
rect 134 1272 137 1278
rect 154 1268 158 1271
rect 202 1268 206 1271
rect 142 1262 145 1268
rect 182 1262 185 1268
rect 238 1262 241 1278
rect 270 1272 273 1278
rect 278 1272 281 1278
rect 318 1272 321 1278
rect 114 1258 118 1261
rect 202 1258 206 1261
rect 158 1252 161 1258
rect 262 1252 265 1258
rect 98 1248 102 1251
rect 130 1248 134 1251
rect 194 1248 201 1251
rect 174 1242 177 1248
rect 122 1238 126 1241
rect 70 1182 73 1218
rect 94 1192 97 1238
rect 174 1192 177 1228
rect 186 1218 190 1221
rect 198 1192 201 1248
rect 226 1238 230 1241
rect 18 1168 22 1171
rect 42 1168 46 1171
rect 122 1168 126 1171
rect 154 1168 158 1171
rect 122 1158 126 1161
rect 22 1142 25 1148
rect 30 1142 33 1158
rect 42 1148 46 1151
rect 54 1132 57 1148
rect 38 1072 41 1078
rect 54 1072 57 1078
rect 62 1062 65 1158
rect 70 1142 73 1148
rect 78 1062 81 1118
rect 86 1092 89 1128
rect 86 1062 89 1068
rect 34 1058 38 1061
rect 62 1052 65 1058
rect 10 1048 14 1051
rect 90 1048 94 1051
rect 22 1042 25 1048
rect 22 992 25 1018
rect 74 988 78 991
rect 86 972 89 1018
rect 102 992 105 1158
rect 110 1152 113 1158
rect 110 1132 113 1148
rect 142 1142 145 1158
rect 166 1152 169 1168
rect 186 1158 193 1161
rect 110 1062 113 1088
rect 126 1082 129 1118
rect 126 1041 129 1078
rect 138 1068 142 1071
rect 150 1052 153 1148
rect 166 1142 169 1148
rect 178 1128 182 1131
rect 190 1122 193 1158
rect 166 1082 169 1088
rect 198 1082 201 1188
rect 206 1162 209 1218
rect 206 1112 209 1138
rect 214 1132 217 1138
rect 162 1068 166 1071
rect 210 1058 214 1061
rect 122 1038 129 1041
rect 18 968 22 971
rect 58 968 62 971
rect 90 958 94 961
rect 6 862 9 938
rect 14 892 17 948
rect 30 942 33 958
rect 66 948 70 951
rect 34 938 38 941
rect 14 872 17 888
rect 6 852 9 858
rect 22 792 25 928
rect 46 922 49 948
rect 38 892 41 918
rect 46 881 49 918
rect 78 892 81 958
rect 126 951 129 1018
rect 142 952 145 1018
rect 174 1011 177 1058
rect 222 1052 225 1158
rect 238 1152 241 1248
rect 250 1238 254 1241
rect 270 1232 273 1268
rect 306 1258 310 1261
rect 294 1232 297 1258
rect 318 1192 321 1268
rect 270 1172 273 1178
rect 254 1162 257 1168
rect 254 1148 262 1151
rect 230 1142 233 1148
rect 230 1102 233 1138
rect 238 1132 241 1138
rect 254 1132 257 1148
rect 286 1142 289 1158
rect 266 1138 273 1141
rect 254 1092 257 1128
rect 270 1112 273 1138
rect 270 1092 273 1108
rect 286 1082 289 1138
rect 294 1132 297 1148
rect 302 1142 305 1158
rect 318 1142 321 1188
rect 342 1182 345 1268
rect 406 1262 409 1278
rect 418 1268 422 1271
rect 458 1268 462 1271
rect 354 1258 358 1261
rect 426 1258 430 1261
rect 366 1242 369 1249
rect 386 1248 390 1251
rect 334 1162 337 1168
rect 358 1162 361 1228
rect 382 1212 385 1238
rect 382 1192 385 1208
rect 370 1168 374 1171
rect 390 1162 393 1178
rect 334 1142 337 1148
rect 302 1122 305 1138
rect 342 1132 345 1148
rect 302 1092 305 1118
rect 318 1112 321 1128
rect 342 1122 345 1128
rect 350 1112 353 1158
rect 362 1148 366 1151
rect 398 1151 401 1258
rect 414 1242 417 1248
rect 406 1192 409 1238
rect 446 1232 449 1248
rect 454 1221 457 1258
rect 478 1242 481 1278
rect 510 1262 513 1268
rect 598 1262 601 1268
rect 614 1262 617 1278
rect 622 1262 625 1278
rect 634 1268 638 1271
rect 650 1268 654 1271
rect 666 1268 670 1271
rect 686 1262 689 1268
rect 718 1262 721 1278
rect 790 1272 793 1278
rect 778 1268 782 1271
rect 742 1262 745 1268
rect 846 1262 849 1268
rect 894 1262 897 1268
rect 810 1258 814 1261
rect 502 1252 505 1258
rect 550 1252 553 1258
rect 514 1238 518 1241
rect 530 1238 542 1241
rect 446 1218 457 1221
rect 446 1192 449 1218
rect 550 1212 553 1218
rect 480 1203 482 1207
rect 486 1203 489 1207
rect 493 1203 496 1207
rect 550 1192 553 1198
rect 558 1192 561 1248
rect 598 1232 601 1258
rect 598 1202 601 1228
rect 590 1182 593 1188
rect 422 1162 425 1178
rect 434 1168 438 1171
rect 398 1148 406 1151
rect 426 1148 430 1151
rect 398 1132 401 1148
rect 410 1138 414 1141
rect 366 1092 369 1128
rect 454 1122 457 1128
rect 430 1092 433 1118
rect 402 1088 406 1091
rect 354 1078 358 1081
rect 246 1072 249 1078
rect 254 1062 257 1078
rect 186 1048 190 1051
rect 202 1038 206 1041
rect 234 1038 238 1041
rect 214 1032 217 1038
rect 246 1032 249 1058
rect 262 1042 265 1078
rect 390 1072 393 1078
rect 462 1072 465 1118
rect 470 1072 473 1138
rect 278 1032 281 1068
rect 166 1008 177 1011
rect 166 992 169 1008
rect 158 962 161 968
rect 166 952 169 968
rect 182 961 185 1018
rect 222 992 225 1028
rect 294 992 297 1048
rect 302 1032 305 1058
rect 322 1048 326 1051
rect 314 1038 318 1041
rect 326 992 329 1038
rect 334 1032 337 1058
rect 342 1042 345 1068
rect 374 1062 377 1068
rect 406 1062 409 1068
rect 426 1058 430 1061
rect 350 1052 353 1058
rect 382 1052 385 1058
rect 406 1042 409 1058
rect 426 1048 430 1051
rect 438 1042 441 1068
rect 458 1058 462 1061
rect 482 1058 486 1061
rect 502 1052 505 1118
rect 510 1082 513 1128
rect 518 1092 521 1138
rect 510 1062 513 1068
rect 534 1062 537 1158
rect 614 1142 617 1148
rect 578 1138 582 1141
rect 602 1138 606 1141
rect 542 1132 545 1138
rect 562 1128 566 1131
rect 622 1131 625 1258
rect 654 1252 657 1258
rect 694 1248 710 1251
rect 738 1248 742 1251
rect 646 1192 649 1198
rect 678 1192 681 1248
rect 694 1242 697 1248
rect 730 1238 734 1241
rect 702 1232 705 1238
rect 742 1192 745 1218
rect 758 1192 761 1258
rect 818 1248 822 1251
rect 718 1172 721 1178
rect 746 1168 750 1171
rect 614 1128 625 1131
rect 674 1158 678 1161
rect 630 1142 633 1158
rect 682 1148 686 1151
rect 662 1142 665 1148
rect 642 1138 646 1141
rect 630 1132 633 1138
rect 662 1132 665 1138
rect 642 1128 646 1131
rect 598 1122 601 1128
rect 550 1062 553 1078
rect 454 992 457 1048
rect 474 1038 478 1041
rect 462 992 465 1028
rect 510 1012 513 1058
rect 518 1032 521 1038
rect 534 1032 537 1048
rect 550 1042 553 1048
rect 558 1022 561 1068
rect 480 1003 482 1007
rect 486 1003 489 1007
rect 493 1003 496 1007
rect 566 992 569 1108
rect 614 1092 617 1128
rect 606 1072 609 1088
rect 622 1082 625 1088
rect 662 1082 665 1088
rect 646 1072 649 1078
rect 586 1068 590 1071
rect 630 1062 633 1068
rect 578 1058 582 1061
rect 590 1042 593 1058
rect 598 1052 601 1058
rect 590 992 593 1008
rect 622 992 625 1038
rect 514 988 518 991
rect 178 958 185 961
rect 182 952 185 958
rect 126 948 137 951
rect 86 932 89 938
rect 74 888 78 891
rect 102 882 105 918
rect 38 878 49 881
rect 30 862 33 878
rect 38 852 41 878
rect 66 868 70 871
rect 50 858 54 861
rect 14 672 17 768
rect 30 762 33 818
rect 38 792 41 848
rect 78 842 81 878
rect 86 862 89 868
rect 98 858 102 861
rect 78 792 81 838
rect 6 652 9 658
rect 6 522 9 528
rect 14 451 17 668
rect 22 652 25 748
rect 30 682 33 758
rect 38 752 41 758
rect 54 752 57 788
rect 66 758 70 761
rect 62 742 65 748
rect 78 742 81 768
rect 86 752 89 838
rect 94 822 97 848
rect 98 758 102 761
rect 98 748 102 751
rect 46 701 49 738
rect 86 732 89 748
rect 98 728 102 731
rect 46 698 57 701
rect 46 682 49 688
rect 54 682 57 698
rect 110 692 113 948
rect 134 942 137 948
rect 190 942 193 968
rect 234 958 238 961
rect 118 932 121 938
rect 126 932 129 938
rect 206 932 209 958
rect 222 942 225 948
rect 262 942 265 978
rect 286 972 289 978
rect 318 972 321 978
rect 382 972 385 978
rect 406 972 409 978
rect 470 972 473 978
rect 518 972 521 978
rect 542 972 545 978
rect 394 968 398 971
rect 434 968 438 971
rect 246 932 249 938
rect 270 932 273 948
rect 254 922 257 928
rect 142 892 145 898
rect 254 892 257 908
rect 218 888 222 891
rect 122 868 126 871
rect 146 858 150 861
rect 126 822 129 858
rect 158 852 161 888
rect 250 868 254 871
rect 174 862 177 868
rect 182 862 185 868
rect 154 848 158 851
rect 158 792 161 838
rect 166 822 169 848
rect 174 812 177 858
rect 198 852 201 868
rect 270 862 273 868
rect 254 852 257 858
rect 186 838 190 841
rect 270 792 273 858
rect 278 852 281 858
rect 286 852 289 858
rect 294 852 297 948
rect 302 932 305 958
rect 322 948 326 951
rect 334 922 337 958
rect 342 932 345 968
rect 406 958 422 961
rect 350 942 353 948
rect 358 942 361 948
rect 366 942 369 948
rect 374 942 377 958
rect 386 948 390 951
rect 406 942 409 958
rect 418 938 422 941
rect 326 918 334 921
rect 302 872 305 878
rect 326 862 329 918
rect 414 892 417 938
rect 366 888 374 891
rect 338 868 342 871
rect 130 758 134 761
rect 126 752 129 758
rect 142 752 145 788
rect 118 732 121 738
rect 126 692 129 748
rect 150 742 153 768
rect 198 762 201 768
rect 170 758 174 761
rect 250 758 254 761
rect 274 758 278 761
rect 202 748 206 751
rect 54 662 57 678
rect 82 668 86 671
rect 86 652 89 658
rect 94 652 97 658
rect 102 652 105 658
rect 54 572 57 578
rect 42 568 46 571
rect 34 548 38 551
rect 22 470 25 478
rect 38 472 41 518
rect 62 492 65 648
rect 70 492 73 538
rect 78 532 81 628
rect 86 572 89 638
rect 102 572 105 648
rect 110 642 113 668
rect 110 561 113 638
rect 118 572 121 648
rect 134 592 137 738
rect 182 732 185 738
rect 142 642 145 658
rect 150 652 153 708
rect 166 692 169 728
rect 162 658 166 661
rect 174 652 177 728
rect 190 662 193 738
rect 214 722 217 758
rect 222 732 225 738
rect 230 692 233 748
rect 270 742 273 748
rect 294 742 297 748
rect 274 728 278 731
rect 254 722 257 728
rect 206 662 209 688
rect 214 672 217 678
rect 222 662 225 688
rect 242 678 246 681
rect 238 662 241 668
rect 254 662 257 718
rect 262 712 265 728
rect 278 672 281 698
rect 302 692 305 858
rect 342 852 345 858
rect 358 852 361 858
rect 366 852 369 888
rect 374 882 377 888
rect 406 872 409 878
rect 430 872 433 948
rect 454 922 457 958
rect 462 952 465 968
rect 502 941 505 958
rect 510 952 513 968
rect 534 942 537 958
rect 542 952 545 958
rect 502 938 513 941
rect 502 932 505 938
rect 438 892 441 918
rect 510 892 513 938
rect 550 922 553 968
rect 446 872 449 888
rect 378 868 382 871
rect 394 868 398 871
rect 482 868 486 871
rect 530 868 534 871
rect 422 862 425 868
rect 394 858 398 861
rect 446 852 449 858
rect 314 848 318 851
rect 434 848 438 851
rect 354 838 358 841
rect 326 832 329 838
rect 406 822 409 848
rect 318 692 321 738
rect 310 682 313 688
rect 286 672 289 678
rect 326 672 329 818
rect 454 782 457 848
rect 430 772 433 778
rect 334 762 337 768
rect 358 762 361 768
rect 334 742 337 748
rect 342 702 345 728
rect 350 722 353 758
rect 358 752 361 758
rect 374 742 377 758
rect 398 742 401 768
rect 406 752 409 758
rect 386 738 390 741
rect 350 702 353 718
rect 342 692 345 698
rect 358 692 361 718
rect 366 692 369 698
rect 306 668 310 671
rect 374 671 377 738
rect 422 732 425 768
rect 438 752 441 758
rect 430 742 433 748
rect 462 742 465 828
rect 470 752 473 858
rect 478 852 481 858
rect 480 803 482 807
rect 486 803 489 807
rect 493 803 496 807
rect 502 792 505 868
rect 526 852 529 858
rect 518 842 521 848
rect 534 842 537 848
rect 494 762 497 778
rect 510 772 513 798
rect 526 772 529 778
rect 502 752 505 768
rect 534 762 537 808
rect 542 801 545 888
rect 566 882 569 948
rect 598 942 601 968
rect 614 951 617 958
rect 614 948 622 951
rect 586 928 593 931
rect 590 892 593 928
rect 586 878 590 881
rect 574 872 577 878
rect 550 812 553 848
rect 558 842 561 858
rect 566 822 569 868
rect 542 798 553 801
rect 550 792 553 798
rect 558 782 561 798
rect 558 772 561 778
rect 458 738 462 741
rect 442 728 446 731
rect 382 702 385 728
rect 454 722 457 728
rect 390 708 398 711
rect 382 682 385 698
rect 390 692 393 708
rect 446 692 449 718
rect 454 682 457 688
rect 470 672 473 748
rect 534 732 537 758
rect 566 752 569 818
rect 574 762 577 838
rect 582 791 585 878
rect 590 832 593 848
rect 598 842 601 938
rect 606 922 609 948
rect 622 932 625 948
rect 630 892 633 1058
rect 638 1052 641 1058
rect 670 1052 673 1148
rect 678 1072 681 1138
rect 694 1132 697 1168
rect 706 1148 710 1151
rect 710 1122 713 1138
rect 690 1068 694 1071
rect 678 1062 681 1068
rect 710 1062 713 1078
rect 718 1072 721 1148
rect 734 1142 737 1158
rect 754 1148 758 1151
rect 766 1092 769 1158
rect 790 1152 793 1198
rect 806 1152 809 1238
rect 814 1182 817 1218
rect 838 1162 841 1188
rect 774 1132 777 1148
rect 806 1092 809 1118
rect 814 1112 817 1158
rect 846 1152 849 1258
rect 862 1231 865 1250
rect 910 1191 913 1278
rect 1102 1272 1105 1278
rect 950 1262 953 1268
rect 1034 1258 1038 1261
rect 994 1218 998 1221
rect 902 1188 913 1191
rect 838 1092 841 1128
rect 886 1111 889 1138
rect 902 1132 905 1188
rect 998 1152 1001 1218
rect 1018 1168 1022 1171
rect 982 1122 985 1128
rect 998 1122 1001 1148
rect 1030 1132 1033 1248
rect 1038 1222 1041 1248
rect 1086 1192 1089 1268
rect 1226 1258 1230 1261
rect 1230 1222 1233 1248
rect 1182 1212 1185 1218
rect 1066 1188 1070 1191
rect 1054 1161 1057 1188
rect 1098 1168 1102 1171
rect 1110 1162 1113 1168
rect 1054 1158 1065 1161
rect 1050 1148 1054 1151
rect 1062 1142 1065 1158
rect 1122 1158 1126 1161
rect 1086 1152 1089 1158
rect 1110 1152 1113 1158
rect 1050 1138 1054 1141
rect 1074 1138 1078 1141
rect 1026 1128 1030 1131
rect 886 1108 897 1111
rect 870 1092 873 1108
rect 894 1092 897 1108
rect 862 1082 865 1088
rect 730 1078 734 1081
rect 906 1078 910 1081
rect 782 1072 785 1078
rect 730 1068 734 1071
rect 762 1068 769 1071
rect 742 1062 745 1068
rect 694 1052 697 1058
rect 650 1048 654 1051
rect 666 1048 670 1051
rect 702 1042 705 1058
rect 750 1052 753 1058
rect 758 1052 761 1058
rect 722 1048 726 1051
rect 654 992 657 1018
rect 694 992 697 1028
rect 706 968 710 971
rect 646 942 649 948
rect 638 932 641 938
rect 646 922 649 938
rect 654 932 657 968
rect 766 962 769 1068
rect 774 982 777 1048
rect 798 1022 801 1078
rect 918 1072 921 1098
rect 926 1092 929 1108
rect 958 1082 961 1118
rect 982 1082 985 1118
rect 1000 1103 1002 1107
rect 1006 1103 1009 1107
rect 1013 1103 1016 1107
rect 998 1082 1001 1088
rect 966 1072 969 1078
rect 882 1068 886 1071
rect 814 1042 817 1068
rect 834 1058 838 1061
rect 914 1058 918 1061
rect 946 1058 950 1061
rect 970 1058 974 1061
rect 822 992 825 1058
rect 830 992 833 1048
rect 838 1022 841 1048
rect 850 1038 854 1041
rect 878 1032 881 1058
rect 858 988 862 991
rect 678 952 681 958
rect 686 941 689 958
rect 682 938 689 941
rect 638 892 641 908
rect 670 892 673 938
rect 614 872 617 878
rect 606 812 609 868
rect 630 862 633 868
rect 614 832 617 848
rect 630 832 633 858
rect 638 852 641 858
rect 582 788 593 791
rect 602 788 606 791
rect 582 772 585 778
rect 590 772 593 788
rect 578 758 582 761
rect 546 748 550 751
rect 578 748 582 751
rect 606 742 609 748
rect 526 692 529 728
rect 534 692 537 728
rect 550 672 553 678
rect 558 672 561 688
rect 574 672 577 708
rect 606 682 609 718
rect 614 692 617 778
rect 630 762 633 798
rect 646 792 649 838
rect 622 732 625 748
rect 598 678 606 681
rect 370 668 377 671
rect 386 668 390 671
rect 194 658 198 661
rect 270 652 273 658
rect 326 652 329 668
rect 334 662 337 668
rect 142 612 145 638
rect 150 562 153 648
rect 158 642 161 648
rect 286 642 289 648
rect 166 631 169 638
rect 158 628 169 631
rect 158 602 161 628
rect 110 558 121 561
rect 78 482 81 528
rect 86 472 89 518
rect 102 492 105 548
rect 110 542 113 548
rect 94 472 97 488
rect 30 452 33 468
rect 54 462 57 468
rect 74 458 78 461
rect 14 448 25 451
rect 58 448 62 451
rect 6 362 9 418
rect 22 392 25 448
rect 78 392 81 438
rect 86 422 89 448
rect 82 368 86 371
rect 70 352 73 358
rect 26 348 30 351
rect 42 348 46 351
rect 82 348 86 351
rect 34 338 38 341
rect 46 312 49 338
rect 54 332 57 338
rect 62 332 65 338
rect 70 331 73 348
rect 78 342 81 348
rect 70 328 81 331
rect 70 292 73 318
rect 6 272 9 288
rect 54 272 57 278
rect 78 262 81 328
rect 94 282 97 468
rect 110 452 113 478
rect 110 392 113 438
rect 118 432 121 558
rect 150 552 153 558
rect 130 548 134 551
rect 134 512 137 548
rect 158 542 161 598
rect 190 592 193 638
rect 258 628 262 631
rect 214 592 217 608
rect 246 582 249 588
rect 198 572 201 578
rect 226 568 230 571
rect 178 558 182 561
rect 190 552 193 558
rect 226 548 230 551
rect 238 542 241 558
rect 146 538 150 541
rect 254 541 257 568
rect 318 562 321 578
rect 274 558 281 561
rect 266 548 273 551
rect 254 538 265 541
rect 174 532 177 538
rect 174 522 177 528
rect 142 462 145 468
rect 158 452 161 518
rect 166 502 169 518
rect 182 482 185 488
rect 166 472 169 478
rect 190 472 193 478
rect 238 472 241 498
rect 246 482 249 538
rect 254 492 257 508
rect 262 472 265 538
rect 270 482 273 548
rect 278 532 281 558
rect 298 548 302 551
rect 310 542 313 558
rect 282 528 286 531
rect 294 522 297 538
rect 282 518 286 521
rect 190 462 193 468
rect 170 458 174 461
rect 142 442 145 448
rect 142 392 145 428
rect 150 372 153 378
rect 126 362 129 368
rect 102 332 105 338
rect 102 272 105 308
rect 110 292 113 348
rect 134 322 137 358
rect 142 322 145 348
rect 158 342 161 448
rect 190 392 193 458
rect 206 392 209 418
rect 214 382 217 418
rect 210 368 214 371
rect 238 371 241 468
rect 270 462 273 478
rect 318 472 321 548
rect 326 522 329 568
rect 334 562 337 658
rect 346 648 350 651
rect 394 648 398 651
rect 366 642 369 648
rect 350 592 353 598
rect 362 568 366 571
rect 306 468 310 471
rect 298 458 302 461
rect 278 442 281 448
rect 230 368 241 371
rect 166 342 169 348
rect 182 342 185 368
rect 150 292 153 338
rect 158 292 161 338
rect 170 328 174 331
rect 182 281 185 338
rect 190 292 193 318
rect 182 278 193 281
rect 74 258 78 261
rect 90 258 94 261
rect 22 192 25 258
rect 82 248 86 251
rect 38 242 41 248
rect 102 242 105 268
rect 118 252 121 278
rect 138 268 142 271
rect 158 242 161 268
rect 166 252 169 258
rect 174 252 177 268
rect 86 192 89 238
rect 182 192 185 258
rect 190 242 193 278
rect 198 262 201 358
rect 230 352 233 368
rect 250 358 254 361
rect 210 348 214 351
rect 206 332 209 348
rect 230 342 233 348
rect 278 342 281 388
rect 286 362 289 448
rect 310 442 313 448
rect 310 392 313 438
rect 286 331 289 358
rect 326 352 329 358
rect 278 328 289 331
rect 206 272 209 278
rect 218 268 222 271
rect 206 262 209 268
rect 222 252 225 258
rect 238 242 241 298
rect 246 252 249 258
rect 254 252 257 258
rect 270 242 273 268
rect 278 262 281 328
rect 302 322 305 338
rect 322 328 326 331
rect 286 302 289 318
rect 302 292 305 318
rect 194 238 198 241
rect 198 182 201 188
rect 246 182 249 218
rect 14 172 17 178
rect 150 172 153 178
rect 22 152 25 158
rect 30 92 33 158
rect 38 152 41 158
rect 46 132 49 168
rect 62 162 65 168
rect 166 162 169 168
rect 74 158 81 161
rect 58 148 62 151
rect 54 72 57 88
rect 62 82 65 138
rect 78 92 81 158
rect 138 158 142 161
rect 94 122 97 138
rect 102 132 105 158
rect 130 148 134 151
rect 118 132 121 138
rect 102 102 105 128
rect 126 92 129 118
rect 62 72 65 78
rect 118 72 121 88
rect 158 62 161 138
rect 166 82 169 158
rect 182 152 185 158
rect 174 112 177 148
rect 190 142 193 158
rect 190 122 193 138
rect 174 72 177 108
rect 206 92 209 168
rect 214 152 217 158
rect 230 152 233 158
rect 238 132 241 148
rect 246 142 249 168
rect 182 72 185 88
rect 230 72 233 98
rect 238 82 241 118
rect 246 92 249 138
rect 254 92 257 238
rect 278 232 281 258
rect 286 252 289 288
rect 298 268 302 271
rect 326 262 329 278
rect 334 262 337 558
rect 342 532 345 558
rect 354 548 358 551
rect 374 542 377 568
rect 398 552 401 648
rect 422 632 425 668
rect 422 552 425 628
rect 430 552 433 658
rect 446 552 449 618
rect 454 592 457 648
rect 480 603 482 607
rect 486 603 489 607
rect 493 603 496 607
rect 502 592 505 668
rect 582 662 585 678
rect 598 672 601 678
rect 490 588 494 591
rect 510 552 513 658
rect 410 548 414 551
rect 374 492 377 518
rect 382 482 385 548
rect 390 542 393 548
rect 426 538 430 541
rect 414 531 417 538
rect 414 528 422 531
rect 438 512 441 538
rect 446 521 449 548
rect 454 532 457 548
rect 462 522 465 528
rect 446 518 457 521
rect 434 478 438 481
rect 358 472 361 478
rect 342 452 345 468
rect 398 462 401 468
rect 406 462 409 478
rect 386 458 390 461
rect 342 392 345 428
rect 350 372 353 458
rect 366 392 369 448
rect 406 442 409 448
rect 422 442 425 478
rect 434 468 438 471
rect 446 451 449 468
rect 454 462 457 518
rect 470 502 473 538
rect 510 532 513 538
rect 526 532 529 648
rect 534 642 537 648
rect 558 592 561 628
rect 566 552 569 658
rect 598 652 601 658
rect 578 588 582 591
rect 598 562 601 648
rect 606 612 609 668
rect 614 592 617 688
rect 630 682 633 758
rect 646 692 649 748
rect 654 712 657 858
rect 662 852 665 868
rect 674 848 681 851
rect 662 752 665 848
rect 670 792 673 838
rect 678 771 681 848
rect 686 842 689 938
rect 694 952 697 958
rect 742 952 745 958
rect 774 952 777 978
rect 870 972 873 1018
rect 786 968 790 971
rect 814 952 817 958
rect 870 952 873 958
rect 754 948 758 951
rect 802 948 806 951
rect 694 912 697 948
rect 718 942 721 948
rect 730 938 734 941
rect 750 932 753 938
rect 722 928 726 931
rect 766 922 769 948
rect 778 938 782 941
rect 678 768 686 771
rect 686 762 689 768
rect 694 751 697 858
rect 702 792 705 868
rect 686 748 697 751
rect 710 752 713 918
rect 718 872 721 908
rect 790 892 793 948
rect 806 922 809 938
rect 814 902 817 948
rect 830 932 833 948
rect 838 922 841 938
rect 838 892 841 918
rect 846 892 849 918
rect 878 892 881 1018
rect 910 992 913 1038
rect 990 1012 993 1078
rect 1038 1062 1041 1138
rect 1134 1132 1137 1208
rect 1166 1192 1169 1198
rect 1198 1162 1201 1218
rect 1210 1158 1214 1161
rect 1142 1152 1145 1158
rect 1246 1152 1249 1258
rect 1278 1202 1281 1268
rect 1294 1221 1297 1278
rect 1454 1272 1457 1278
rect 1430 1262 1433 1268
rect 1406 1232 1409 1238
rect 1414 1222 1417 1258
rect 1438 1252 1441 1258
rect 1294 1218 1305 1221
rect 1254 1160 1257 1188
rect 1218 1148 1225 1151
rect 1166 1142 1169 1148
rect 1174 1142 1177 1148
rect 1146 1138 1150 1141
rect 1182 1132 1185 1148
rect 1206 1142 1209 1148
rect 1194 1138 1198 1141
rect 1110 1102 1113 1118
rect 1110 1082 1113 1088
rect 1210 1078 1214 1081
rect 894 962 897 978
rect 966 972 969 978
rect 954 968 958 971
rect 974 962 977 988
rect 990 962 993 968
rect 1022 962 1025 1058
rect 1062 1031 1065 1050
rect 1062 992 1065 1008
rect 1094 992 1097 1068
rect 1150 1042 1153 1058
rect 1202 1048 1206 1051
rect 1158 992 1161 1048
rect 1194 1018 1198 1021
rect 1202 988 1206 991
rect 1054 962 1057 978
rect 966 952 969 958
rect 922 948 926 951
rect 886 902 889 938
rect 910 922 913 948
rect 922 938 926 941
rect 938 928 942 931
rect 926 901 929 928
rect 918 898 929 901
rect 738 888 742 891
rect 870 882 873 888
rect 918 882 921 898
rect 930 888 934 891
rect 946 878 950 881
rect 862 872 865 878
rect 746 868 750 871
rect 758 862 761 868
rect 726 802 729 848
rect 734 822 737 848
rect 758 812 761 858
rect 722 788 726 791
rect 662 692 665 738
rect 686 722 689 748
rect 694 722 697 728
rect 710 692 713 748
rect 726 742 729 748
rect 718 722 721 738
rect 682 688 686 691
rect 710 682 713 688
rect 642 678 646 681
rect 698 678 702 681
rect 674 668 678 671
rect 622 602 625 668
rect 634 658 638 661
rect 638 592 641 628
rect 618 558 622 561
rect 538 548 542 551
rect 602 548 606 551
rect 538 538 542 541
rect 566 531 569 548
rect 566 528 574 531
rect 518 522 521 528
rect 498 478 502 481
rect 462 472 465 478
rect 490 468 494 471
rect 478 462 481 468
rect 510 462 513 478
rect 518 472 521 508
rect 534 492 537 528
rect 550 522 553 528
rect 550 502 553 518
rect 542 472 545 498
rect 574 492 577 528
rect 590 512 593 538
rect 606 532 609 538
rect 614 492 617 498
rect 578 468 582 471
rect 610 468 614 471
rect 458 458 462 461
rect 446 448 457 451
rect 398 382 401 388
rect 418 368 422 371
rect 350 272 353 368
rect 454 362 457 448
rect 358 322 361 358
rect 382 352 385 358
rect 374 342 377 348
rect 426 338 430 341
rect 366 262 369 328
rect 382 262 385 288
rect 390 272 393 278
rect 278 162 281 218
rect 326 202 329 258
rect 342 242 345 248
rect 406 242 409 288
rect 438 262 441 338
rect 446 302 449 348
rect 454 342 457 358
rect 462 342 465 448
rect 480 403 482 407
rect 486 403 489 407
rect 493 403 496 407
rect 478 342 481 348
rect 446 262 449 298
rect 454 292 457 318
rect 470 272 473 338
rect 462 262 465 268
rect 370 218 374 221
rect 310 162 313 178
rect 290 148 294 151
rect 318 142 321 158
rect 326 152 329 178
rect 342 172 345 178
rect 398 172 401 218
rect 362 168 366 171
rect 350 152 353 158
rect 366 152 369 158
rect 298 138 302 141
rect 374 141 377 158
rect 398 142 401 168
rect 406 152 409 158
rect 414 152 417 258
rect 422 252 425 258
rect 438 252 441 258
rect 430 242 433 248
rect 430 152 433 198
rect 438 162 441 218
rect 446 172 449 238
rect 480 203 482 207
rect 486 203 489 207
rect 493 203 496 207
rect 478 152 481 188
rect 486 152 489 158
rect 502 152 505 258
rect 510 232 513 458
rect 518 452 521 468
rect 526 452 529 458
rect 534 452 537 458
rect 526 432 529 448
rect 550 432 553 468
rect 558 452 561 468
rect 574 452 577 458
rect 518 292 521 398
rect 526 342 529 348
rect 550 342 553 428
rect 558 392 561 448
rect 574 421 577 448
rect 566 418 577 421
rect 558 342 561 348
rect 566 322 569 418
rect 582 412 585 448
rect 574 372 577 378
rect 590 352 593 468
rect 622 462 625 558
rect 630 542 633 578
rect 598 402 601 458
rect 614 442 617 448
rect 622 412 625 418
rect 598 372 601 398
rect 614 392 617 398
rect 526 272 529 318
rect 590 292 593 348
rect 510 152 513 228
rect 374 138 382 141
rect 410 138 414 141
rect 262 132 265 138
rect 278 132 281 138
rect 382 132 385 138
rect 270 62 273 118
rect 302 102 305 118
rect 390 112 393 118
rect 278 72 281 78
rect 286 72 289 98
rect 334 72 337 88
rect 350 82 353 98
rect 358 72 361 108
rect 374 72 377 78
rect 414 72 417 128
rect 154 58 158 61
rect 370 58 374 61
rect 398 52 401 58
rect 258 48 262 51
rect 306 48 310 51
rect 270 -18 273 8
rect 430 -18 433 148
rect 478 142 481 148
rect 510 142 513 148
rect 518 142 521 248
rect 534 242 537 268
rect 566 262 569 268
rect 554 248 558 251
rect 458 138 462 141
rect 518 132 521 138
rect 534 132 537 168
rect 558 162 561 168
rect 546 148 550 151
rect 462 122 465 128
rect 470 72 473 118
rect 494 92 497 128
rect 450 68 454 71
rect 494 62 497 68
rect 482 58 486 61
rect 518 42 521 78
rect 526 62 529 118
rect 534 112 537 128
rect 566 72 569 218
rect 574 72 577 288
rect 598 271 601 348
rect 622 282 625 298
rect 630 292 633 498
rect 638 472 641 518
rect 646 492 649 548
rect 654 482 657 668
rect 662 652 665 658
rect 670 562 673 658
rect 702 652 705 668
rect 670 552 673 558
rect 686 552 689 638
rect 718 582 721 648
rect 726 632 729 738
rect 734 692 737 808
rect 742 762 745 778
rect 750 752 753 798
rect 774 792 777 798
rect 806 782 809 868
rect 818 858 822 861
rect 854 842 857 868
rect 870 852 873 878
rect 914 868 918 871
rect 842 818 846 821
rect 762 768 766 771
rect 750 742 753 748
rect 782 741 785 758
rect 806 742 809 748
rect 814 742 817 798
rect 822 782 825 788
rect 826 758 830 761
rect 858 758 862 761
rect 830 752 833 758
rect 782 738 790 741
rect 750 672 753 688
rect 738 668 742 671
rect 766 661 769 738
rect 782 662 785 718
rect 790 672 793 738
rect 814 732 817 738
rect 830 722 833 738
rect 838 732 841 738
rect 790 662 793 668
rect 766 658 774 661
rect 730 548 734 551
rect 670 532 673 538
rect 678 492 681 518
rect 662 452 665 458
rect 670 352 673 458
rect 686 442 689 548
rect 710 532 713 538
rect 694 492 697 528
rect 702 492 705 508
rect 694 482 697 488
rect 718 472 721 508
rect 726 472 729 478
rect 742 472 745 658
rect 750 612 753 658
rect 766 632 769 658
rect 782 651 785 658
rect 778 648 785 651
rect 766 622 769 628
rect 798 622 801 718
rect 846 692 849 758
rect 862 722 865 748
rect 870 742 873 828
rect 878 792 881 818
rect 886 772 889 868
rect 894 862 897 868
rect 910 832 913 848
rect 934 832 937 868
rect 942 782 945 878
rect 966 862 969 938
rect 966 822 969 858
rect 894 742 897 778
rect 918 762 921 768
rect 942 762 945 778
rect 958 772 961 818
rect 902 742 905 748
rect 950 742 953 758
rect 870 692 873 708
rect 822 672 825 688
rect 814 642 817 658
rect 750 562 753 608
rect 758 562 761 618
rect 806 582 809 618
rect 790 572 793 578
rect 822 572 825 668
rect 854 662 857 668
rect 878 662 881 678
rect 846 602 849 648
rect 810 558 814 561
rect 750 532 753 558
rect 766 532 769 538
rect 762 518 766 521
rect 774 492 777 558
rect 854 551 857 658
rect 846 548 857 551
rect 862 648 870 651
rect 862 552 865 648
rect 878 642 881 658
rect 886 652 889 728
rect 918 722 921 728
rect 894 662 897 678
rect 902 662 905 678
rect 926 662 929 738
rect 942 732 945 738
rect 958 731 961 748
rect 950 728 961 731
rect 950 722 953 728
rect 958 692 961 718
rect 946 678 950 681
rect 966 681 969 818
rect 974 762 977 958
rect 982 922 985 938
rect 990 932 993 948
rect 958 678 969 681
rect 914 658 918 661
rect 902 642 905 648
rect 926 632 929 658
rect 942 652 945 668
rect 930 618 934 621
rect 874 558 878 561
rect 790 512 793 548
rect 798 542 801 548
rect 698 468 702 471
rect 714 468 718 471
rect 750 471 753 478
rect 746 468 753 471
rect 686 352 689 418
rect 702 402 705 448
rect 710 362 713 418
rect 718 352 721 388
rect 690 348 694 351
rect 706 348 710 351
rect 646 322 649 348
rect 694 342 697 348
rect 658 328 662 331
rect 646 282 649 298
rect 654 272 657 288
rect 686 282 689 338
rect 718 332 721 338
rect 726 312 729 448
rect 734 362 737 418
rect 742 392 745 448
rect 750 352 753 468
rect 762 458 766 461
rect 758 392 761 448
rect 774 422 777 468
rect 790 462 793 468
rect 782 452 785 458
rect 766 402 769 418
rect 774 372 777 408
rect 798 392 801 478
rect 822 472 825 488
rect 810 468 814 471
rect 830 462 833 548
rect 846 532 849 548
rect 854 522 857 538
rect 838 512 841 518
rect 862 482 865 548
rect 878 532 881 558
rect 910 552 913 598
rect 926 562 929 568
rect 958 562 961 678
rect 966 662 969 668
rect 974 662 977 748
rect 982 712 985 918
rect 1000 903 1002 907
rect 1006 903 1009 907
rect 1013 903 1016 907
rect 1022 892 1025 958
rect 1074 948 1078 951
rect 1038 942 1041 948
rect 1054 942 1057 948
rect 1030 932 1033 938
rect 1062 882 1065 888
rect 1058 868 1062 871
rect 1038 792 1041 848
rect 1062 842 1065 848
rect 990 742 993 748
rect 1014 732 1017 748
rect 990 691 993 718
rect 1000 703 1002 707
rect 1006 703 1009 707
rect 1013 703 1016 707
rect 990 688 1001 691
rect 982 672 985 678
rect 990 652 993 678
rect 938 548 942 551
rect 886 542 889 548
rect 898 538 902 541
rect 934 532 937 538
rect 894 481 897 518
rect 926 482 929 518
rect 894 478 905 481
rect 878 472 881 478
rect 902 472 905 478
rect 890 468 894 471
rect 930 468 934 471
rect 814 442 817 458
rect 814 432 817 438
rect 754 348 758 351
rect 798 342 801 348
rect 806 342 809 368
rect 822 352 825 358
rect 830 352 833 448
rect 838 372 841 468
rect 950 462 953 538
rect 958 502 961 558
rect 982 552 985 558
rect 970 548 974 551
rect 914 458 918 461
rect 846 382 849 458
rect 854 452 857 458
rect 862 452 865 458
rect 870 432 873 448
rect 854 392 857 428
rect 886 422 889 458
rect 950 452 953 458
rect 958 452 961 468
rect 974 462 977 498
rect 990 492 993 648
rect 998 632 1001 688
rect 1014 602 1017 668
rect 1022 662 1025 788
rect 1062 752 1065 838
rect 1070 792 1073 948
rect 1102 942 1105 948
rect 1142 932 1145 938
rect 1122 928 1129 931
rect 1094 922 1097 928
rect 1094 902 1097 918
rect 1126 892 1129 928
rect 1158 922 1161 948
rect 1174 912 1177 958
rect 1182 942 1185 948
rect 1194 938 1198 941
rect 1214 932 1217 1018
rect 1222 942 1225 1148
rect 1234 1068 1238 1071
rect 1246 1062 1249 1148
rect 1286 1142 1289 1158
rect 1302 1132 1305 1218
rect 1406 1152 1409 1208
rect 1430 1182 1433 1188
rect 1462 1172 1465 1268
rect 1478 1242 1481 1248
rect 1486 1231 1489 1298
rect 1478 1228 1489 1231
rect 1502 1271 1505 1318
rect 1498 1268 1505 1271
rect 1394 1138 1398 1141
rect 1406 1132 1409 1138
rect 1438 1132 1441 1148
rect 1454 1142 1457 1148
rect 1410 1128 1414 1131
rect 1302 1092 1305 1128
rect 1398 1122 1401 1128
rect 1318 1082 1321 1088
rect 1302 1072 1305 1078
rect 1230 952 1233 1058
rect 1246 1042 1249 1058
rect 1254 1022 1257 1048
rect 1254 962 1257 988
rect 1270 952 1273 1058
rect 1218 928 1222 931
rect 1230 912 1233 948
rect 1246 892 1249 918
rect 1198 882 1201 888
rect 1178 878 1182 881
rect 1098 868 1102 871
rect 1162 868 1166 871
rect 1078 802 1081 868
rect 1110 862 1113 868
rect 1118 841 1121 868
rect 1190 862 1193 878
rect 1238 872 1241 878
rect 1226 868 1230 871
rect 1170 858 1174 861
rect 1110 838 1121 841
rect 1142 842 1145 848
rect 1090 818 1094 821
rect 1110 792 1113 838
rect 1078 752 1081 768
rect 1086 752 1089 758
rect 1030 712 1033 738
rect 1054 732 1057 748
rect 1046 681 1049 728
rect 1054 692 1057 718
rect 1046 678 1057 681
rect 1042 668 1046 671
rect 1046 652 1049 658
rect 1006 542 1009 578
rect 1014 562 1017 568
rect 1014 542 1017 548
rect 1038 542 1041 648
rect 1054 582 1057 678
rect 1062 671 1065 718
rect 1070 712 1073 738
rect 1062 668 1073 671
rect 1062 652 1065 658
rect 1070 652 1073 668
rect 1086 662 1089 738
rect 1114 728 1118 731
rect 1118 722 1121 728
rect 1102 671 1105 718
rect 1098 668 1105 671
rect 1110 651 1113 708
rect 1118 662 1121 678
rect 1126 672 1129 808
rect 1190 792 1193 798
rect 1206 772 1209 868
rect 1214 762 1217 768
rect 1134 742 1137 748
rect 1142 742 1145 758
rect 1150 732 1153 748
rect 1190 742 1193 748
rect 1166 702 1169 728
rect 1198 722 1201 748
rect 1222 742 1225 788
rect 1230 742 1233 858
rect 1142 698 1150 701
rect 1142 692 1145 698
rect 1154 678 1158 681
rect 1174 672 1177 678
rect 1106 648 1113 651
rect 1126 652 1129 658
rect 1054 552 1057 578
rect 1062 552 1065 648
rect 1086 562 1089 618
rect 1102 552 1105 558
rect 1050 538 1054 541
rect 1034 528 1038 531
rect 1070 531 1073 548
rect 1110 542 1113 568
rect 1118 552 1121 608
rect 1150 572 1153 668
rect 1162 658 1166 661
rect 1182 652 1185 678
rect 1190 662 1193 678
rect 1206 672 1209 728
rect 1214 672 1217 738
rect 1226 728 1230 731
rect 1238 722 1241 818
rect 1246 742 1249 878
rect 1254 872 1257 878
rect 1262 872 1265 878
rect 1278 862 1281 868
rect 1286 862 1289 898
rect 1302 892 1305 938
rect 1318 932 1321 1078
rect 1398 1052 1401 1118
rect 1454 1081 1457 1098
rect 1462 1091 1465 1148
rect 1470 1112 1473 1218
rect 1478 1192 1481 1228
rect 1462 1088 1470 1091
rect 1454 1078 1462 1081
rect 1414 1062 1417 1068
rect 1462 1062 1465 1068
rect 1418 1058 1422 1061
rect 1434 1058 1438 1061
rect 1474 1058 1478 1061
rect 1426 1048 1430 1051
rect 1399 952 1402 958
rect 1406 952 1409 1038
rect 1446 992 1449 1038
rect 1434 968 1438 971
rect 1478 962 1481 968
rect 1486 952 1489 1218
rect 1494 1202 1497 1268
rect 1466 948 1470 951
rect 1398 892 1401 938
rect 1438 932 1441 948
rect 1454 941 1457 948
rect 1454 938 1465 941
rect 1454 932 1457 938
rect 1410 888 1414 891
rect 1310 872 1313 878
rect 1322 868 1326 871
rect 1266 858 1270 861
rect 1286 832 1289 848
rect 1270 752 1273 788
rect 1286 772 1289 778
rect 1294 762 1297 868
rect 1302 762 1305 858
rect 1358 852 1361 858
rect 1374 852 1377 868
rect 1390 862 1393 868
rect 1318 792 1321 848
rect 1382 842 1385 858
rect 1294 752 1297 758
rect 1254 742 1257 748
rect 1298 738 1302 741
rect 1262 722 1265 738
rect 1238 682 1241 718
rect 1226 678 1230 681
rect 1262 672 1265 678
rect 1270 672 1273 678
rect 1286 672 1289 688
rect 1234 668 1238 671
rect 1206 662 1209 668
rect 1254 662 1257 668
rect 1274 658 1278 661
rect 1242 648 1246 651
rect 1166 592 1169 648
rect 1230 622 1233 648
rect 1254 642 1257 658
rect 1286 652 1289 668
rect 1134 562 1137 568
rect 1206 562 1209 618
rect 1186 558 1190 561
rect 1222 552 1225 558
rect 1162 548 1166 551
rect 1210 548 1214 551
rect 1234 548 1238 551
rect 1246 542 1249 578
rect 1278 552 1281 648
rect 1294 562 1297 698
rect 1302 692 1305 708
rect 1310 682 1313 788
rect 1326 762 1329 768
rect 1318 742 1321 758
rect 1342 752 1345 768
rect 1358 762 1361 798
rect 1358 742 1361 748
rect 1366 742 1369 778
rect 1374 772 1377 778
rect 1398 762 1401 858
rect 1374 752 1377 758
rect 1390 752 1393 758
rect 1330 738 1334 741
rect 1318 672 1321 678
rect 1334 672 1337 688
rect 1366 681 1369 738
rect 1366 678 1377 681
rect 1374 672 1377 678
rect 1326 662 1329 668
rect 1350 662 1353 668
rect 1366 662 1369 668
rect 1302 652 1305 658
rect 1326 642 1329 658
rect 1302 562 1305 568
rect 1294 552 1297 558
rect 1326 552 1329 578
rect 1334 552 1337 558
rect 1342 552 1345 658
rect 1358 651 1361 658
rect 1358 648 1369 651
rect 1358 592 1361 618
rect 1350 572 1353 578
rect 1366 542 1369 648
rect 1374 642 1377 648
rect 1382 562 1385 748
rect 1398 702 1401 758
rect 1406 702 1409 878
rect 1422 862 1425 908
rect 1438 882 1441 928
rect 1450 878 1454 881
rect 1462 862 1465 938
rect 1426 858 1430 861
rect 1486 852 1489 928
rect 1414 792 1417 848
rect 1478 842 1481 848
rect 1462 792 1465 838
rect 1486 822 1489 848
rect 1494 831 1497 918
rect 1502 842 1505 868
rect 1494 828 1505 831
rect 1454 752 1457 758
rect 1414 732 1417 748
rect 1422 742 1425 748
rect 1434 738 1438 741
rect 1430 692 1433 728
rect 1438 692 1441 698
rect 1462 692 1465 718
rect 1470 712 1473 738
rect 1390 672 1393 678
rect 1382 542 1385 558
rect 1090 538 1094 541
rect 1266 538 1270 541
rect 1370 538 1374 541
rect 1070 528 1078 531
rect 1000 503 1002 507
rect 1006 503 1009 507
rect 1013 503 1016 507
rect 1046 492 1049 528
rect 1054 492 1057 528
rect 1078 522 1081 528
rect 990 478 1017 481
rect 990 472 993 478
rect 1014 472 1017 478
rect 1038 472 1041 478
rect 1002 468 1006 471
rect 1026 458 1030 461
rect 938 448 942 451
rect 838 352 841 358
rect 846 352 849 358
rect 814 342 817 348
rect 862 342 865 388
rect 882 368 886 371
rect 750 332 753 338
rect 742 322 745 328
rect 782 312 785 318
rect 738 288 742 291
rect 586 268 601 271
rect 582 232 585 258
rect 590 252 593 258
rect 598 192 601 268
rect 606 192 609 258
rect 614 152 617 268
rect 678 262 681 278
rect 694 272 697 288
rect 710 282 713 288
rect 666 258 670 261
rect 686 252 689 268
rect 634 248 638 251
rect 646 248 654 251
rect 638 152 641 158
rect 582 132 585 148
rect 582 92 585 98
rect 538 68 542 71
rect 562 68 566 71
rect 480 3 482 7
rect 486 3 489 7
rect 493 3 496 7
rect 518 -18 521 38
rect 542 -18 545 58
rect 574 -18 577 68
rect 598 62 601 148
rect 606 82 609 148
rect 614 92 617 148
rect 622 132 625 138
rect 638 92 641 128
rect 646 112 649 248
rect 654 132 657 238
rect 678 152 681 158
rect 702 152 705 278
rect 750 262 753 308
rect 794 288 798 291
rect 774 271 777 288
rect 782 282 785 288
rect 806 282 809 338
rect 790 271 793 278
rect 774 268 793 271
rect 814 272 817 298
rect 822 292 825 338
rect 830 282 833 338
rect 870 332 873 358
rect 902 352 905 358
rect 918 352 921 388
rect 926 352 929 358
rect 886 342 889 348
rect 910 342 913 348
rect 842 328 846 331
rect 890 328 894 331
rect 870 302 873 328
rect 862 282 865 288
rect 838 272 841 278
rect 878 272 881 318
rect 918 282 921 338
rect 942 332 945 378
rect 958 352 961 368
rect 966 341 969 428
rect 974 362 977 458
rect 990 452 993 458
rect 998 452 1001 458
rect 1014 452 1017 458
rect 1054 452 1057 488
rect 1078 472 1081 478
rect 1086 472 1089 518
rect 1066 468 1070 471
rect 1046 432 1049 448
rect 1062 442 1065 458
rect 1086 452 1089 458
rect 1014 352 1017 368
rect 958 338 969 341
rect 1022 342 1025 418
rect 1086 402 1089 418
rect 1050 378 1054 381
rect 1082 378 1086 381
rect 1046 362 1049 368
rect 1030 352 1033 358
rect 1046 342 1049 348
rect 1062 342 1065 368
rect 1074 358 1078 361
rect 1086 341 1089 358
rect 1094 352 1097 528
rect 1134 492 1137 508
rect 1118 482 1121 488
rect 1102 452 1105 468
rect 1102 352 1105 378
rect 1110 362 1113 418
rect 1126 392 1129 478
rect 1150 472 1153 518
rect 1150 462 1153 468
rect 1158 462 1161 538
rect 1190 532 1193 538
rect 1178 468 1182 471
rect 1190 462 1193 528
rect 1158 452 1161 458
rect 1198 451 1201 518
rect 1230 492 1233 528
rect 1254 522 1257 528
rect 1262 511 1265 528
rect 1254 508 1265 511
rect 1210 468 1214 471
rect 1254 471 1257 508
rect 1262 482 1265 488
rect 1254 468 1262 471
rect 1218 458 1222 461
rect 1230 452 1233 468
rect 1246 462 1249 468
rect 1270 462 1273 488
rect 1294 472 1297 518
rect 1318 472 1321 538
rect 1370 518 1374 521
rect 1382 492 1385 498
rect 1346 478 1350 481
rect 1390 481 1393 548
rect 1382 478 1393 481
rect 1398 482 1401 658
rect 1406 642 1409 648
rect 1414 542 1417 658
rect 1422 632 1425 638
rect 1454 622 1457 668
rect 1470 642 1473 678
rect 1486 672 1489 718
rect 1494 662 1497 818
rect 1502 762 1505 828
rect 1442 588 1446 591
rect 1450 548 1454 551
rect 1466 548 1470 551
rect 1498 548 1502 551
rect 1426 538 1430 541
rect 1462 532 1465 538
rect 1486 532 1489 538
rect 1422 522 1425 528
rect 1414 492 1417 508
rect 1346 468 1350 471
rect 1282 458 1286 461
rect 1198 448 1206 451
rect 1174 432 1177 448
rect 1134 352 1137 398
rect 1158 352 1161 418
rect 1174 372 1177 428
rect 1214 402 1217 448
rect 1230 442 1233 448
rect 1238 412 1241 458
rect 1270 442 1273 448
rect 1174 358 1182 361
rect 1118 342 1121 348
rect 1086 338 1094 341
rect 1150 341 1153 348
rect 1150 338 1158 341
rect 958 292 961 338
rect 1114 328 1118 331
rect 982 322 985 328
rect 974 282 977 318
rect 990 302 993 318
rect 1000 303 1002 307
rect 1006 303 1009 307
rect 1013 303 1016 307
rect 1038 292 1041 298
rect 1110 292 1113 318
rect 1126 302 1129 338
rect 1150 292 1153 318
rect 1174 292 1177 358
rect 1194 348 1198 351
rect 1182 322 1185 328
rect 1190 302 1193 338
rect 1206 312 1209 358
rect 1242 348 1246 351
rect 1214 312 1217 328
rect 1222 302 1225 338
rect 1270 332 1273 408
rect 1286 382 1289 388
rect 1294 332 1297 468
rect 1302 452 1305 458
rect 1310 432 1313 458
rect 1318 452 1321 468
rect 1366 462 1369 468
rect 1366 442 1369 448
rect 1382 422 1385 478
rect 1398 472 1401 478
rect 1398 452 1401 458
rect 1142 282 1145 288
rect 962 278 966 281
rect 1154 278 1158 281
rect 1174 278 1182 281
rect 758 262 761 268
rect 894 262 897 268
rect 918 262 921 278
rect 926 262 929 268
rect 842 258 846 261
rect 934 261 937 278
rect 1054 272 1057 278
rect 1102 272 1105 278
rect 1118 272 1121 278
rect 946 268 950 271
rect 978 268 982 271
rect 1002 268 1006 271
rect 934 258 942 261
rect 710 252 713 258
rect 766 252 769 258
rect 742 182 745 188
rect 726 162 729 178
rect 746 168 750 171
rect 750 152 753 158
rect 666 148 670 151
rect 694 142 697 148
rect 702 142 705 148
rect 726 142 729 148
rect 662 121 665 138
rect 654 118 665 121
rect 646 92 649 108
rect 654 82 657 118
rect 662 92 665 98
rect 650 78 654 81
rect 670 62 673 138
rect 734 132 737 148
rect 678 72 681 128
rect 690 118 694 121
rect 714 88 718 91
rect 758 82 761 248
rect 806 232 809 258
rect 858 248 862 251
rect 806 222 809 228
rect 774 202 777 218
rect 798 192 801 208
rect 770 158 774 161
rect 858 158 862 161
rect 802 148 806 151
rect 766 132 769 138
rect 778 128 782 131
rect 698 78 702 81
rect 734 72 737 78
rect 758 72 761 78
rect 682 68 686 71
rect 674 58 681 61
rect 590 22 593 38
rect 598 12 601 58
rect 642 48 646 51
rect 662 42 665 48
rect 638 -18 641 8
rect 662 -18 665 38
rect 678 -18 681 58
rect 686 12 689 68
rect 706 58 710 61
rect 726 52 729 68
rect 738 58 742 61
rect 750 52 753 58
rect 702 -18 705 8
rect 750 -18 753 48
rect 774 -9 777 128
rect 782 82 785 88
rect 794 68 798 71
rect 794 58 798 61
rect 786 48 790 51
rect 794 48 798 51
rect 774 -12 785 -9
rect 782 -18 785 -12
rect 806 -18 809 148
rect 822 92 825 132
rect 854 112 857 138
rect 862 132 865 148
rect 830 92 833 108
rect 862 92 865 118
rect 870 92 873 248
rect 930 238 937 241
rect 878 152 881 158
rect 886 142 889 218
rect 934 192 937 238
rect 942 232 945 258
rect 990 252 993 258
rect 942 162 945 178
rect 958 152 961 168
rect 902 142 905 148
rect 910 142 913 148
rect 894 112 897 138
rect 918 132 921 138
rect 814 52 817 88
rect 822 62 825 78
rect 846 72 849 78
rect 862 72 865 78
rect 910 72 913 78
rect 942 72 945 128
rect 962 88 966 91
rect 982 72 985 178
rect 1014 152 1017 268
rect 1026 266 1030 269
rect 1054 252 1057 268
rect 1078 262 1081 268
rect 1074 248 1078 251
rect 1046 222 1049 238
rect 1042 218 1046 221
rect 990 142 993 148
rect 922 68 926 71
rect 846 62 849 68
rect 902 62 905 68
rect 950 62 953 68
rect 990 62 993 138
rect 998 132 1001 138
rect 1000 103 1002 107
rect 1006 103 1009 107
rect 1013 103 1016 107
rect 1006 72 1009 78
rect 1022 72 1025 128
rect 1038 81 1041 198
rect 1070 172 1073 228
rect 1086 202 1089 268
rect 1094 252 1097 258
rect 1126 222 1129 258
rect 1134 242 1137 268
rect 1158 262 1161 268
rect 1166 262 1169 268
rect 1174 261 1177 278
rect 1214 272 1217 288
rect 1270 282 1273 328
rect 1286 272 1289 298
rect 1186 268 1190 271
rect 1242 268 1246 271
rect 1298 268 1302 271
rect 1310 271 1313 418
rect 1334 412 1337 418
rect 1406 412 1409 468
rect 1334 392 1337 398
rect 1358 372 1361 408
rect 1366 392 1369 408
rect 1414 392 1417 428
rect 1378 358 1382 361
rect 1362 348 1366 351
rect 1378 348 1382 351
rect 1342 342 1345 348
rect 1318 322 1321 338
rect 1330 328 1334 331
rect 1310 268 1321 271
rect 1174 258 1185 261
rect 1242 258 1246 261
rect 1274 258 1278 261
rect 1058 168 1062 171
rect 1046 158 1070 161
rect 1046 152 1049 158
rect 1102 152 1105 158
rect 1118 152 1121 208
rect 1134 162 1137 198
rect 1134 152 1137 158
rect 1054 142 1057 148
rect 1046 132 1049 138
rect 1070 92 1073 148
rect 1142 142 1145 178
rect 1154 168 1158 171
rect 1098 138 1102 141
rect 1078 122 1081 138
rect 1110 132 1113 138
rect 1078 102 1081 118
rect 1094 92 1097 128
rect 1118 122 1121 128
rect 1038 78 1046 81
rect 930 58 934 61
rect 938 58 945 61
rect 1018 58 1022 61
rect 1034 58 1038 61
rect 1070 61 1073 88
rect 1102 62 1105 108
rect 1110 82 1113 98
rect 1126 82 1129 128
rect 1150 102 1153 148
rect 1182 141 1185 258
rect 1194 248 1198 251
rect 1222 232 1225 248
rect 1262 222 1265 258
rect 1230 192 1233 198
rect 1198 151 1201 168
rect 1194 148 1201 151
rect 1214 151 1217 158
rect 1210 148 1217 151
rect 1182 138 1193 141
rect 1166 92 1169 128
rect 1174 112 1177 118
rect 1190 92 1193 138
rect 1206 122 1209 138
rect 1246 132 1249 208
rect 1262 192 1265 218
rect 1286 212 1289 268
rect 1306 258 1310 261
rect 1262 142 1265 168
rect 1270 152 1273 188
rect 1282 168 1286 171
rect 1318 162 1321 268
rect 1326 262 1329 278
rect 1334 262 1337 268
rect 1326 192 1329 258
rect 1334 172 1337 188
rect 1342 182 1345 338
rect 1382 292 1385 328
rect 1390 282 1393 358
rect 1410 348 1414 351
rect 1402 338 1406 341
rect 1414 332 1417 348
rect 1422 342 1425 518
rect 1430 452 1433 528
rect 1478 502 1481 528
rect 1486 482 1489 518
rect 1494 511 1497 518
rect 1494 508 1502 511
rect 1494 492 1497 498
rect 1478 472 1481 478
rect 1454 452 1457 458
rect 1486 372 1489 478
rect 1502 462 1505 488
rect 1438 362 1441 368
rect 1434 348 1438 351
rect 1486 342 1489 368
rect 1434 328 1438 331
rect 1402 288 1406 291
rect 1438 282 1441 328
rect 1454 322 1457 338
rect 1370 268 1374 271
rect 1390 262 1393 278
rect 1418 268 1422 271
rect 1358 172 1361 248
rect 1306 158 1310 161
rect 1386 158 1390 161
rect 1366 152 1369 158
rect 1278 148 1286 151
rect 1338 148 1350 151
rect 1126 72 1129 78
rect 1066 58 1073 61
rect 1114 58 1118 61
rect 1142 61 1145 88
rect 1278 82 1281 148
rect 1354 138 1361 141
rect 1370 138 1374 141
rect 1286 132 1289 138
rect 1358 132 1361 138
rect 1346 128 1350 131
rect 1310 122 1313 128
rect 1154 78 1166 81
rect 1234 78 1238 81
rect 1222 72 1225 78
rect 1246 72 1249 78
rect 1294 72 1297 88
rect 1342 82 1345 88
rect 1366 72 1369 78
rect 1374 72 1377 118
rect 1382 92 1385 148
rect 1398 122 1401 148
rect 1406 142 1409 178
rect 1414 121 1417 258
rect 1430 232 1433 268
rect 1438 262 1441 278
rect 1454 272 1457 278
rect 1462 262 1465 318
rect 1478 282 1481 338
rect 1486 322 1489 328
rect 1486 282 1489 318
rect 1502 292 1505 458
rect 1462 192 1465 248
rect 1478 152 1481 158
rect 1442 148 1449 151
rect 1490 148 1494 151
rect 1422 132 1425 138
rect 1414 118 1425 121
rect 1414 92 1417 108
rect 1422 82 1425 118
rect 1430 112 1433 128
rect 1446 92 1449 148
rect 1438 72 1441 78
rect 1454 72 1457 78
rect 1462 72 1465 78
rect 1154 68 1158 71
rect 1178 68 1182 71
rect 1234 68 1238 71
rect 1290 68 1294 71
rect 1330 68 1337 71
rect 1482 68 1486 71
rect 1198 62 1201 68
rect 1142 58 1150 61
rect 1210 58 1214 61
rect 862 52 865 58
rect 886 52 889 58
rect 942 51 945 58
rect 958 51 961 58
rect 1078 52 1081 58
rect 942 48 961 51
rect 1026 48 1030 51
rect 1194 48 1198 51
rect 1206 -18 1209 48
rect 1246 42 1249 68
rect 1298 58 1302 61
rect 1322 58 1326 61
rect 1254 22 1257 58
rect 1334 52 1337 68
rect 1374 62 1377 68
rect 1426 58 1430 61
rect 1466 58 1470 61
rect 1398 52 1401 58
rect 1494 52 1497 148
rect 1502 132 1505 258
rect 1314 48 1318 51
rect 1270 21 1273 48
rect 1266 18 1273 21
rect 1262 -18 1265 18
rect 270 -22 274 -18
rect 430 -22 434 -18
rect 518 -22 522 -18
rect 542 -22 546 -18
rect 574 -22 578 -18
rect 638 -22 642 -18
rect 662 -22 666 -18
rect 678 -22 682 -18
rect 702 -22 706 -18
rect 750 -22 754 -18
rect 782 -22 786 -18
rect 806 -22 810 -18
rect 1206 -22 1210 -18
rect 1262 -22 1266 -18
<< m3contact >>
rect 102 1288 106 1292
rect 462 1288 466 1292
rect 70 1278 74 1282
rect 6 1268 10 1272
rect 14 1268 18 1272
rect 38 1268 42 1272
rect 22 1238 26 1242
rect 38 1238 42 1242
rect 94 1258 98 1262
rect 1518 1318 1522 1322
rect 1002 1303 1006 1307
rect 1009 1303 1013 1307
rect 1486 1298 1490 1302
rect 134 1278 138 1282
rect 238 1278 242 1282
rect 270 1278 274 1282
rect 278 1278 282 1282
rect 406 1278 410 1282
rect 566 1278 570 1282
rect 622 1278 626 1282
rect 654 1278 658 1282
rect 774 1278 778 1282
rect 790 1278 794 1282
rect 910 1278 914 1282
rect 1214 1278 1218 1282
rect 1374 1278 1378 1282
rect 142 1268 146 1272
rect 150 1268 154 1272
rect 182 1268 186 1272
rect 206 1268 210 1272
rect 318 1268 322 1272
rect 118 1258 122 1262
rect 158 1258 162 1262
rect 206 1258 210 1262
rect 86 1248 90 1252
rect 94 1248 98 1252
rect 134 1248 138 1252
rect 174 1248 178 1252
rect 94 1238 98 1242
rect 126 1238 130 1242
rect 30 1208 34 1212
rect 62 1208 66 1212
rect 174 1228 178 1232
rect 190 1218 194 1222
rect 238 1248 242 1252
rect 262 1248 266 1252
rect 230 1238 234 1242
rect 198 1188 202 1192
rect 70 1178 74 1182
rect 22 1168 26 1172
rect 38 1168 42 1172
rect 118 1168 122 1172
rect 150 1168 154 1172
rect 166 1168 170 1172
rect 62 1158 66 1162
rect 110 1158 114 1162
rect 126 1158 130 1162
rect 142 1158 146 1162
rect 46 1148 50 1152
rect 22 1138 26 1142
rect 30 1138 34 1142
rect 54 1128 58 1132
rect 54 1078 58 1082
rect 38 1068 42 1072
rect 70 1148 74 1152
rect 86 1088 90 1092
rect 86 1068 90 1072
rect 38 1058 42 1062
rect 78 1058 82 1062
rect 14 1048 18 1052
rect 22 1048 26 1052
rect 62 1048 66 1052
rect 86 1048 90 1052
rect 22 1018 26 1022
rect 78 988 82 992
rect 150 1148 154 1152
rect 110 1128 114 1132
rect 110 1088 114 1092
rect 126 1078 130 1082
rect 142 1068 146 1072
rect 166 1138 170 1142
rect 174 1128 178 1132
rect 190 1118 194 1122
rect 206 1158 210 1162
rect 222 1158 226 1162
rect 214 1128 218 1132
rect 206 1108 210 1112
rect 166 1078 170 1082
rect 198 1078 202 1082
rect 166 1068 170 1072
rect 174 1058 178 1062
rect 206 1058 210 1062
rect 150 1048 154 1052
rect 102 988 106 992
rect 22 968 26 972
rect 54 968 58 972
rect 86 968 90 972
rect 94 958 98 962
rect 6 938 10 942
rect 46 948 50 952
rect 62 948 66 952
rect 30 938 34 942
rect 22 928 26 932
rect 14 888 18 892
rect 6 848 10 852
rect 38 918 42 922
rect 254 1238 258 1242
rect 310 1258 314 1262
rect 270 1228 274 1232
rect 294 1228 298 1232
rect 270 1178 274 1182
rect 254 1158 258 1162
rect 302 1158 306 1162
rect 238 1148 242 1152
rect 238 1128 242 1132
rect 230 1098 234 1102
rect 286 1138 290 1142
rect 270 1108 274 1112
rect 254 1088 258 1092
rect 414 1268 418 1272
rect 454 1268 458 1272
rect 358 1258 362 1262
rect 398 1258 402 1262
rect 422 1258 426 1262
rect 454 1258 458 1262
rect 382 1248 386 1252
rect 366 1238 370 1242
rect 382 1238 386 1242
rect 358 1228 362 1232
rect 342 1178 346 1182
rect 382 1208 386 1212
rect 390 1178 394 1182
rect 366 1168 370 1172
rect 334 1158 338 1162
rect 334 1148 338 1152
rect 318 1138 322 1142
rect 294 1128 298 1132
rect 342 1128 346 1132
rect 302 1118 306 1122
rect 342 1118 346 1122
rect 358 1148 362 1152
rect 414 1238 418 1242
rect 446 1228 450 1232
rect 510 1268 514 1272
rect 598 1268 602 1272
rect 638 1268 642 1272
rect 646 1268 650 1272
rect 670 1268 674 1272
rect 686 1268 690 1272
rect 742 1268 746 1272
rect 774 1268 778 1272
rect 846 1268 850 1272
rect 502 1258 506 1262
rect 614 1258 618 1262
rect 654 1258 658 1262
rect 718 1258 722 1262
rect 758 1258 762 1262
rect 806 1258 810 1262
rect 894 1258 898 1262
rect 550 1248 554 1252
rect 558 1248 562 1252
rect 478 1238 482 1242
rect 510 1238 514 1242
rect 550 1208 554 1212
rect 482 1203 486 1207
rect 489 1203 493 1207
rect 550 1198 554 1202
rect 598 1228 602 1232
rect 598 1198 602 1202
rect 558 1188 562 1192
rect 422 1178 426 1182
rect 590 1178 594 1182
rect 430 1168 434 1172
rect 422 1148 426 1152
rect 406 1138 410 1142
rect 366 1128 370 1132
rect 398 1128 402 1132
rect 318 1108 322 1112
rect 350 1108 354 1112
rect 430 1118 434 1122
rect 454 1118 458 1122
rect 406 1088 410 1092
rect 254 1078 258 1082
rect 286 1078 290 1082
rect 350 1078 354 1082
rect 246 1068 250 1072
rect 182 1048 186 1052
rect 198 1038 202 1042
rect 214 1038 218 1042
rect 230 1038 234 1042
rect 342 1068 346 1072
rect 390 1068 394 1072
rect 438 1068 442 1072
rect 462 1068 466 1072
rect 470 1068 474 1072
rect 262 1038 266 1042
rect 294 1048 298 1052
rect 222 1028 226 1032
rect 246 1028 250 1032
rect 278 1028 282 1032
rect 166 968 170 972
rect 158 958 162 962
rect 318 1048 322 1052
rect 318 1038 322 1042
rect 326 1038 330 1042
rect 302 1028 306 1032
rect 350 1058 354 1062
rect 374 1058 378 1062
rect 406 1058 410 1062
rect 422 1058 426 1062
rect 382 1048 386 1052
rect 430 1048 434 1052
rect 454 1058 458 1062
rect 478 1058 482 1062
rect 518 1088 522 1092
rect 510 1078 514 1082
rect 510 1068 514 1072
rect 614 1148 618 1152
rect 582 1138 586 1142
rect 606 1138 610 1142
rect 542 1128 546 1132
rect 558 1128 562 1132
rect 734 1248 738 1252
rect 646 1198 650 1202
rect 726 1238 730 1242
rect 702 1228 706 1232
rect 814 1248 818 1252
rect 790 1198 794 1202
rect 678 1188 682 1192
rect 742 1188 746 1192
rect 718 1178 722 1182
rect 742 1168 746 1172
rect 630 1158 634 1162
rect 670 1158 674 1162
rect 662 1148 666 1152
rect 670 1148 674 1152
rect 678 1148 682 1152
rect 630 1138 634 1142
rect 646 1138 650 1142
rect 638 1128 642 1132
rect 662 1128 666 1132
rect 598 1118 602 1122
rect 566 1108 570 1112
rect 550 1078 554 1082
rect 558 1068 562 1072
rect 534 1058 538 1062
rect 454 1048 458 1052
rect 406 1038 410 1042
rect 334 1028 338 1032
rect 478 1038 482 1042
rect 462 1028 466 1032
rect 550 1048 554 1052
rect 518 1028 522 1032
rect 534 1028 538 1032
rect 558 1018 562 1022
rect 510 1008 514 1012
rect 482 1003 486 1007
rect 489 1003 493 1007
rect 606 1088 610 1092
rect 622 1088 626 1092
rect 646 1078 650 1082
rect 662 1078 666 1082
rect 582 1068 586 1072
rect 582 1058 586 1062
rect 630 1058 634 1062
rect 598 1048 602 1052
rect 590 1038 594 1042
rect 622 1038 626 1042
rect 590 1008 594 1012
rect 454 988 458 992
rect 518 988 522 992
rect 262 978 266 982
rect 286 978 290 982
rect 318 978 322 982
rect 382 978 386 982
rect 406 978 410 982
rect 470 978 474 982
rect 518 978 522 982
rect 190 968 194 972
rect 86 928 90 932
rect 102 918 106 922
rect 70 888 74 892
rect 78 878 82 882
rect 102 878 106 882
rect 30 858 34 862
rect 70 868 74 872
rect 46 858 50 862
rect 86 868 90 872
rect 94 858 98 862
rect 86 838 90 842
rect 38 788 42 792
rect 54 788 58 792
rect 78 788 82 792
rect 38 758 42 762
rect 6 648 10 652
rect 6 518 10 522
rect 62 758 66 762
rect 62 748 66 752
rect 94 818 98 822
rect 102 758 106 762
rect 94 748 98 752
rect 78 738 82 742
rect 86 728 90 732
rect 94 728 98 732
rect 206 958 210 962
rect 230 958 234 962
rect 342 968 346 972
rect 398 968 402 972
rect 430 968 434 972
rect 462 968 466 972
rect 510 968 514 972
rect 542 968 546 972
rect 294 948 298 952
rect 222 938 226 942
rect 246 938 250 942
rect 118 928 122 932
rect 126 928 130 932
rect 254 928 258 932
rect 270 928 274 932
rect 254 908 258 912
rect 142 898 146 902
rect 158 888 162 892
rect 214 888 218 892
rect 126 868 130 872
rect 142 858 146 862
rect 174 868 178 872
rect 254 868 258 872
rect 270 868 274 872
rect 182 858 186 862
rect 150 848 154 852
rect 126 818 130 822
rect 166 818 170 822
rect 278 858 282 862
rect 198 848 202 852
rect 254 848 258 852
rect 190 838 194 842
rect 174 808 178 812
rect 318 948 322 952
rect 302 928 306 932
rect 374 958 378 962
rect 350 948 354 952
rect 358 948 362 952
rect 390 948 394 952
rect 366 938 370 942
rect 374 938 378 942
rect 406 938 410 942
rect 422 938 426 942
rect 334 918 338 922
rect 302 878 306 882
rect 374 888 378 892
rect 414 888 418 892
rect 342 868 346 872
rect 342 858 346 862
rect 286 848 290 852
rect 294 848 298 852
rect 142 788 146 792
rect 270 788 274 792
rect 126 758 130 762
rect 198 768 202 772
rect 118 728 122 732
rect 174 758 178 762
rect 254 758 258 762
rect 270 758 274 762
rect 206 748 210 752
rect 134 738 138 742
rect 150 738 154 742
rect 190 738 194 742
rect 46 678 50 682
rect 86 668 90 672
rect 110 668 114 672
rect 54 658 58 662
rect 94 658 98 662
rect 22 648 26 652
rect 62 648 66 652
rect 86 648 90 652
rect 102 648 106 652
rect 54 578 58 582
rect 46 568 50 572
rect 38 548 42 552
rect 22 478 26 482
rect 86 638 90 642
rect 78 628 82 632
rect 118 648 122 652
rect 102 568 106 572
rect 166 728 170 732
rect 182 728 186 732
rect 150 708 154 712
rect 142 658 146 662
rect 158 658 162 662
rect 230 748 234 752
rect 270 748 274 752
rect 222 728 226 732
rect 214 718 218 722
rect 294 738 298 742
rect 254 728 258 732
rect 270 728 274 732
rect 254 718 258 722
rect 206 688 210 692
rect 222 688 226 692
rect 214 678 218 682
rect 246 678 250 682
rect 262 708 266 712
rect 278 698 282 702
rect 406 878 410 882
rect 542 958 546 962
rect 534 938 538 942
rect 502 928 506 932
rect 438 918 442 922
rect 454 918 458 922
rect 550 918 554 922
rect 446 888 450 892
rect 542 888 546 892
rect 382 868 386 872
rect 398 868 402 872
rect 430 868 434 872
rect 486 868 490 872
rect 534 868 538 872
rect 390 858 394 862
rect 422 858 426 862
rect 470 858 474 862
rect 318 848 322 852
rect 358 848 362 852
rect 438 848 442 852
rect 446 848 450 852
rect 358 838 362 842
rect 326 828 330 832
rect 326 818 330 822
rect 406 818 410 822
rect 302 688 306 692
rect 310 688 314 692
rect 286 678 290 682
rect 462 828 466 832
rect 454 778 458 782
rect 334 768 338 772
rect 358 768 362 772
rect 398 768 402 772
rect 430 768 434 772
rect 374 758 378 762
rect 334 738 338 742
rect 342 728 346 732
rect 358 748 362 752
rect 406 758 410 762
rect 390 738 394 742
rect 398 738 402 742
rect 350 718 354 722
rect 342 698 346 702
rect 350 698 354 702
rect 366 698 370 702
rect 358 688 362 692
rect 310 668 314 672
rect 334 668 338 672
rect 366 668 370 672
rect 438 748 442 752
rect 478 848 482 852
rect 482 803 486 807
rect 489 803 493 807
rect 526 848 530 852
rect 534 848 538 852
rect 518 838 522 842
rect 534 808 538 812
rect 510 798 514 802
rect 494 778 498 782
rect 502 768 506 772
rect 526 768 530 772
rect 622 948 626 952
rect 598 938 602 942
rect 566 878 570 882
rect 574 878 578 882
rect 590 878 594 882
rect 558 838 562 842
rect 574 838 578 842
rect 566 818 570 822
rect 550 808 554 812
rect 558 798 562 802
rect 558 778 562 782
rect 470 748 474 752
rect 502 748 506 752
rect 430 738 434 742
rect 454 738 458 742
rect 422 728 426 732
rect 438 728 442 732
rect 446 718 450 722
rect 454 718 458 722
rect 398 708 402 712
rect 382 698 386 702
rect 382 678 386 682
rect 454 678 458 682
rect 606 918 610 922
rect 678 1138 682 1142
rect 702 1148 706 1152
rect 694 1128 698 1132
rect 710 1118 714 1122
rect 710 1078 714 1082
rect 678 1068 682 1072
rect 694 1068 698 1072
rect 750 1148 754 1152
rect 734 1138 738 1142
rect 814 1178 818 1182
rect 774 1148 778 1152
rect 806 1118 810 1122
rect 1102 1268 1106 1272
rect 950 1258 954 1262
rect 1030 1258 1034 1262
rect 1030 1248 1034 1252
rect 998 1218 1002 1222
rect 838 1128 842 1132
rect 814 1108 818 1112
rect 870 1108 874 1112
rect 1014 1168 1018 1172
rect 982 1128 986 1132
rect 1222 1258 1226 1262
rect 1134 1208 1138 1212
rect 1182 1208 1186 1212
rect 1054 1188 1058 1192
rect 1070 1188 1074 1192
rect 1086 1188 1090 1192
rect 1094 1168 1098 1172
rect 1046 1148 1050 1152
rect 1086 1158 1090 1162
rect 1110 1158 1114 1162
rect 1126 1158 1130 1162
rect 1046 1138 1050 1142
rect 1070 1138 1074 1142
rect 1022 1128 1026 1132
rect 958 1118 962 1122
rect 998 1118 1002 1122
rect 926 1108 930 1112
rect 918 1098 922 1102
rect 766 1088 770 1092
rect 862 1088 866 1092
rect 734 1078 738 1082
rect 910 1078 914 1082
rect 718 1068 722 1072
rect 734 1068 738 1072
rect 782 1068 786 1072
rect 694 1058 698 1062
rect 702 1058 706 1062
rect 742 1058 746 1062
rect 758 1058 762 1062
rect 638 1048 642 1052
rect 646 1048 650 1052
rect 670 1048 674 1052
rect 726 1048 730 1052
rect 750 1048 754 1052
rect 694 1028 698 1032
rect 654 1018 658 1022
rect 654 968 658 972
rect 710 968 714 972
rect 646 938 650 942
rect 638 928 642 932
rect 1002 1103 1006 1107
rect 1009 1103 1013 1107
rect 966 1078 970 1082
rect 998 1078 1002 1082
rect 878 1068 882 1072
rect 822 1058 826 1062
rect 830 1058 834 1062
rect 918 1058 922 1062
rect 950 1058 954 1062
rect 974 1058 978 1062
rect 814 1038 818 1042
rect 798 1018 802 1022
rect 830 1048 834 1052
rect 854 1038 858 1042
rect 910 1038 914 1042
rect 878 1028 882 1032
rect 838 1018 842 1022
rect 878 1018 882 1022
rect 822 988 826 992
rect 862 988 866 992
rect 774 978 778 982
rect 678 958 682 962
rect 694 958 698 962
rect 742 958 746 962
rect 766 958 770 962
rect 670 938 674 942
rect 646 918 650 922
rect 638 908 642 912
rect 630 888 634 892
rect 614 878 618 882
rect 606 868 610 872
rect 598 838 602 842
rect 590 828 594 832
rect 630 858 634 862
rect 638 858 642 862
rect 646 838 650 842
rect 614 828 618 832
rect 630 828 634 832
rect 606 808 610 812
rect 630 798 634 802
rect 598 788 602 792
rect 614 778 618 782
rect 582 768 586 772
rect 582 758 586 762
rect 542 748 546 752
rect 566 748 570 752
rect 574 748 578 752
rect 606 738 610 742
rect 526 728 530 732
rect 606 718 610 722
rect 574 708 578 712
rect 558 688 562 692
rect 550 678 554 682
rect 622 748 626 752
rect 614 688 618 692
rect 582 678 586 682
rect 390 668 394 672
rect 470 668 474 672
rect 198 658 202 662
rect 238 658 242 662
rect 174 648 178 652
rect 270 648 274 652
rect 326 648 330 652
rect 142 638 146 642
rect 142 608 146 612
rect 158 638 162 642
rect 190 638 194 642
rect 286 638 290 642
rect 158 598 162 602
rect 102 548 106 552
rect 110 548 114 552
rect 70 488 74 492
rect 78 478 82 482
rect 94 488 98 492
rect 110 478 114 482
rect 38 468 42 472
rect 86 468 90 472
rect 54 458 58 462
rect 70 458 74 462
rect 30 448 34 452
rect 62 448 66 452
rect 86 418 90 422
rect 78 368 82 372
rect 30 348 34 352
rect 46 348 50 352
rect 70 348 74 352
rect 86 348 90 352
rect 38 338 42 342
rect 62 338 66 342
rect 54 328 58 332
rect 78 338 82 342
rect 70 318 74 322
rect 46 308 50 312
rect 6 288 10 292
rect 54 278 58 282
rect 110 438 114 442
rect 150 558 154 562
rect 126 548 130 552
rect 262 628 266 632
rect 214 608 218 612
rect 246 588 250 592
rect 198 578 202 582
rect 230 568 234 572
rect 254 568 258 572
rect 174 558 178 562
rect 190 558 194 562
rect 222 548 226 552
rect 150 538 154 542
rect 174 538 178 542
rect 238 538 242 542
rect 246 538 250 542
rect 326 568 330 572
rect 262 548 266 552
rect 158 518 162 522
rect 174 518 178 522
rect 134 508 138 512
rect 142 468 146 472
rect 166 498 170 502
rect 238 498 242 502
rect 182 488 186 492
rect 190 478 194 482
rect 254 508 258 512
rect 318 558 322 562
rect 294 548 298 552
rect 318 548 322 552
rect 310 538 314 542
rect 286 528 290 532
rect 278 518 282 522
rect 294 518 298 522
rect 270 478 274 482
rect 166 468 170 472
rect 174 458 178 462
rect 190 458 194 462
rect 142 438 146 442
rect 118 428 122 432
rect 142 428 146 432
rect 150 378 154 382
rect 126 368 130 372
rect 102 328 106 332
rect 102 308 106 312
rect 94 278 98 282
rect 206 418 210 422
rect 190 388 194 392
rect 214 378 218 382
rect 182 368 186 372
rect 206 368 210 372
rect 350 648 354 652
rect 398 648 402 652
rect 366 638 370 642
rect 350 598 354 602
rect 366 568 370 572
rect 374 568 378 572
rect 334 558 338 562
rect 326 518 330 522
rect 310 468 314 472
rect 302 458 306 462
rect 286 448 290 452
rect 278 438 282 442
rect 278 388 282 392
rect 166 348 170 352
rect 150 338 154 342
rect 158 338 162 342
rect 134 318 138 322
rect 142 318 146 322
rect 174 328 178 332
rect 158 288 162 292
rect 190 318 194 322
rect 22 258 26 262
rect 70 258 74 262
rect 86 258 90 262
rect 38 248 42 252
rect 78 248 82 252
rect 134 268 138 272
rect 174 268 178 272
rect 118 248 122 252
rect 182 258 186 262
rect 166 248 170 252
rect 86 238 90 242
rect 102 238 106 242
rect 158 238 162 242
rect 254 358 258 362
rect 214 348 218 352
rect 230 348 234 352
rect 310 438 314 442
rect 326 358 330 362
rect 206 328 210 332
rect 238 298 242 302
rect 206 278 210 282
rect 214 268 218 272
rect 198 258 202 262
rect 206 258 210 262
rect 222 248 226 252
rect 270 268 274 272
rect 254 258 258 262
rect 246 248 250 252
rect 326 328 330 332
rect 302 318 306 322
rect 286 298 290 302
rect 286 288 290 292
rect 302 288 306 292
rect 198 238 202 242
rect 254 238 258 242
rect 182 188 186 192
rect 14 178 18 182
rect 198 178 202 182
rect 246 178 250 182
rect 62 168 66 172
rect 150 168 154 172
rect 166 168 170 172
rect 22 158 26 162
rect 38 158 42 162
rect 62 148 66 152
rect 62 138 66 142
rect 46 128 50 132
rect 54 88 58 92
rect 30 78 34 82
rect 102 158 106 162
rect 142 158 146 162
rect 166 158 170 162
rect 182 158 186 162
rect 134 148 138 152
rect 118 128 122 132
rect 94 118 98 122
rect 126 118 130 122
rect 102 98 106 102
rect 118 88 122 92
rect 62 78 66 82
rect 190 138 194 142
rect 190 118 194 122
rect 174 108 178 112
rect 214 158 218 162
rect 230 148 234 152
rect 246 138 250 142
rect 238 128 242 132
rect 238 118 242 122
rect 230 98 234 102
rect 182 88 186 92
rect 326 278 330 282
rect 302 268 306 272
rect 358 548 362 552
rect 422 628 426 632
rect 446 618 450 622
rect 482 603 486 607
rect 489 603 493 607
rect 454 588 458 592
rect 486 588 490 592
rect 502 588 506 592
rect 526 648 530 652
rect 390 548 394 552
rect 406 548 410 552
rect 422 548 426 552
rect 454 548 458 552
rect 342 528 346 532
rect 374 518 378 522
rect 430 538 434 542
rect 462 518 466 522
rect 438 508 442 512
rect 358 478 362 482
rect 382 478 386 482
rect 406 478 410 482
rect 438 478 442 482
rect 382 458 386 462
rect 398 458 402 462
rect 342 448 346 452
rect 342 428 346 432
rect 406 448 410 452
rect 438 468 442 472
rect 534 638 538 642
rect 558 628 562 632
rect 598 648 602 652
rect 582 588 586 592
rect 606 608 610 612
rect 662 848 666 852
rect 670 838 674 842
rect 790 968 794 972
rect 870 968 874 972
rect 870 958 874 962
rect 718 948 722 952
rect 758 948 762 952
rect 766 948 770 952
rect 774 948 778 952
rect 790 948 794 952
rect 806 948 810 952
rect 814 948 818 952
rect 726 938 730 942
rect 726 928 730 932
rect 750 928 754 932
rect 782 938 786 942
rect 710 918 714 922
rect 766 918 770 922
rect 694 908 698 912
rect 686 838 690 842
rect 686 768 690 772
rect 662 748 666 752
rect 718 908 722 912
rect 806 918 810 922
rect 830 928 834 932
rect 838 918 842 922
rect 846 918 850 922
rect 814 898 818 902
rect 1166 1198 1170 1202
rect 1142 1158 1146 1162
rect 1198 1158 1202 1162
rect 1214 1158 1218 1162
rect 1454 1268 1458 1272
rect 1430 1258 1434 1262
rect 1406 1238 1410 1242
rect 1438 1248 1442 1252
rect 1414 1218 1418 1222
rect 1278 1198 1282 1202
rect 1286 1158 1290 1162
rect 1166 1148 1170 1152
rect 1174 1148 1178 1152
rect 1206 1148 1210 1152
rect 1142 1138 1146 1142
rect 1198 1138 1202 1142
rect 1182 1128 1186 1132
rect 1110 1098 1114 1102
rect 1110 1088 1114 1092
rect 1214 1078 1218 1082
rect 1038 1058 1042 1062
rect 990 1008 994 1012
rect 974 988 978 992
rect 894 978 898 982
rect 966 978 970 982
rect 950 968 954 972
rect 990 968 994 972
rect 1062 1008 1066 1012
rect 1158 1048 1162 1052
rect 1198 1048 1202 1052
rect 1150 1038 1154 1042
rect 1198 1018 1202 1022
rect 1214 1018 1218 1022
rect 1094 988 1098 992
rect 1198 988 1202 992
rect 1054 978 1058 982
rect 966 958 970 962
rect 918 948 922 952
rect 926 938 930 942
rect 966 938 970 942
rect 934 928 938 932
rect 910 918 914 922
rect 886 898 890 902
rect 742 888 746 892
rect 870 888 874 892
rect 878 888 882 892
rect 934 888 938 892
rect 862 878 866 882
rect 942 878 946 882
rect 742 868 746 872
rect 758 858 762 862
rect 734 818 738 822
rect 734 808 738 812
rect 758 808 762 812
rect 726 798 730 802
rect 718 788 722 792
rect 654 708 658 712
rect 686 718 690 722
rect 694 718 698 722
rect 726 738 730 742
rect 718 718 722 722
rect 662 688 666 692
rect 678 688 682 692
rect 630 678 634 682
rect 646 678 650 682
rect 702 678 706 682
rect 710 678 714 682
rect 622 668 626 672
rect 670 668 674 672
rect 638 658 642 662
rect 638 628 642 632
rect 622 598 626 602
rect 630 578 634 582
rect 598 558 602 562
rect 614 558 618 562
rect 534 548 538 552
rect 606 548 610 552
rect 542 538 546 542
rect 510 528 514 532
rect 526 528 530 532
rect 534 528 538 532
rect 518 518 522 522
rect 518 508 522 512
rect 470 498 474 502
rect 462 478 466 482
rect 494 478 498 482
rect 510 478 514 482
rect 486 468 490 472
rect 550 518 554 522
rect 542 498 546 502
rect 550 498 554 502
rect 606 528 610 532
rect 590 508 594 512
rect 614 498 618 502
rect 542 468 546 472
rect 582 468 586 472
rect 590 468 594 472
rect 614 468 618 472
rect 462 458 466 462
rect 478 458 482 462
rect 510 458 514 462
rect 422 438 426 442
rect 398 378 402 382
rect 350 368 354 372
rect 414 368 418 372
rect 462 448 466 452
rect 382 358 386 362
rect 374 348 378 352
rect 430 338 434 342
rect 366 328 370 332
rect 358 318 362 322
rect 382 288 386 292
rect 406 288 410 292
rect 390 278 394 282
rect 334 258 338 262
rect 278 228 282 232
rect 482 403 486 407
rect 489 403 493 407
rect 478 348 482 352
rect 462 338 466 342
rect 446 298 450 302
rect 454 288 458 292
rect 470 268 474 272
rect 422 258 426 262
rect 446 258 450 262
rect 462 258 466 262
rect 342 238 346 242
rect 374 218 378 222
rect 326 198 330 202
rect 310 178 314 182
rect 326 178 330 182
rect 342 178 346 182
rect 278 158 282 162
rect 318 158 322 162
rect 294 148 298 152
rect 366 168 370 172
rect 398 168 402 172
rect 350 158 354 162
rect 366 158 370 162
rect 262 138 266 142
rect 302 138 306 142
rect 318 138 322 142
rect 406 158 410 162
rect 438 248 442 252
rect 430 238 434 242
rect 430 198 434 202
rect 482 203 486 207
rect 489 203 493 207
rect 478 188 482 192
rect 446 168 450 172
rect 438 158 442 162
rect 486 158 490 162
rect 534 458 538 462
rect 518 448 522 452
rect 526 448 530 452
rect 574 458 578 462
rect 558 448 562 452
rect 526 428 530 432
rect 550 428 554 432
rect 518 398 522 402
rect 558 388 562 392
rect 526 338 530 342
rect 558 338 562 342
rect 582 408 586 412
rect 574 368 578 372
rect 646 548 650 552
rect 630 498 634 502
rect 622 458 626 462
rect 614 438 618 442
rect 622 408 626 412
rect 598 398 602 402
rect 614 398 618 402
rect 598 368 602 372
rect 526 318 530 322
rect 566 318 570 322
rect 574 288 578 292
rect 590 288 594 292
rect 566 268 570 272
rect 518 248 522 252
rect 510 228 514 232
rect 414 148 418 152
rect 478 148 482 152
rect 502 148 506 152
rect 382 138 386 142
rect 406 138 410 142
rect 278 128 282 132
rect 358 108 362 112
rect 390 108 394 112
rect 286 98 290 102
rect 302 98 306 102
rect 350 98 354 102
rect 278 78 282 82
rect 334 88 338 92
rect 374 78 378 82
rect 414 68 418 72
rect 158 58 162 62
rect 374 58 378 62
rect 398 58 402 62
rect 262 48 266 52
rect 310 48 314 52
rect 270 8 274 12
rect 558 248 562 252
rect 534 238 538 242
rect 566 218 570 222
rect 534 168 538 172
rect 558 168 562 172
rect 462 138 466 142
rect 510 138 514 142
rect 550 148 554 152
rect 494 128 498 132
rect 518 128 522 132
rect 462 118 466 122
rect 518 78 522 82
rect 454 68 458 72
rect 494 68 498 72
rect 486 58 490 62
rect 534 108 538 112
rect 622 298 626 302
rect 662 648 666 652
rect 702 648 706 652
rect 686 638 690 642
rect 670 558 674 562
rect 750 798 754 802
rect 774 798 778 802
rect 742 778 746 782
rect 814 858 818 862
rect 894 868 898 872
rect 910 868 914 872
rect 870 848 874 852
rect 854 838 858 842
rect 870 828 874 832
rect 838 818 842 822
rect 814 798 818 802
rect 806 778 810 782
rect 758 768 762 772
rect 782 758 786 762
rect 750 748 754 752
rect 806 748 810 752
rect 822 778 826 782
rect 822 758 826 762
rect 846 758 850 762
rect 854 758 858 762
rect 830 748 834 752
rect 750 688 754 692
rect 734 668 738 672
rect 742 658 746 662
rect 814 728 818 732
rect 838 728 842 732
rect 798 718 802 722
rect 830 718 834 722
rect 790 668 794 672
rect 782 658 786 662
rect 726 628 730 632
rect 718 578 722 582
rect 670 548 674 552
rect 726 548 730 552
rect 670 538 674 542
rect 678 488 682 492
rect 654 478 658 482
rect 638 468 642 472
rect 670 458 674 462
rect 662 448 666 452
rect 710 538 714 542
rect 702 508 706 512
rect 718 508 722 512
rect 694 488 698 492
rect 694 478 698 482
rect 726 478 730 482
rect 766 628 770 632
rect 878 818 882 822
rect 910 828 914 832
rect 934 828 938 832
rect 958 818 962 822
rect 966 818 970 822
rect 894 778 898 782
rect 942 778 946 782
rect 886 768 890 772
rect 918 768 922 772
rect 958 768 962 772
rect 950 758 954 762
rect 902 738 906 742
rect 918 728 922 732
rect 862 718 866 722
rect 870 708 874 712
rect 822 688 826 692
rect 814 638 818 642
rect 766 618 770 622
rect 798 618 802 622
rect 750 608 754 612
rect 790 578 794 582
rect 806 578 810 582
rect 854 658 858 662
rect 878 658 882 662
rect 846 598 850 602
rect 750 558 754 562
rect 758 558 762 562
rect 814 558 818 562
rect 766 528 770 532
rect 766 518 770 522
rect 798 548 802 552
rect 894 678 898 682
rect 942 728 946 732
rect 950 718 954 722
rect 958 718 962 722
rect 942 678 946 682
rect 990 948 994 952
rect 990 928 994 932
rect 982 918 986 922
rect 974 758 978 762
rect 974 748 978 752
rect 942 668 946 672
rect 902 658 906 662
rect 910 658 914 662
rect 886 648 890 652
rect 878 638 882 642
rect 902 638 906 642
rect 926 628 930 632
rect 934 618 938 622
rect 910 598 914 602
rect 870 558 874 562
rect 790 508 794 512
rect 774 488 778 492
rect 822 488 826 492
rect 750 478 754 482
rect 694 468 698 472
rect 710 468 714 472
rect 686 438 690 442
rect 702 398 706 402
rect 718 388 722 392
rect 710 348 714 352
rect 694 338 698 342
rect 654 328 658 332
rect 646 318 650 322
rect 646 298 650 302
rect 654 288 658 292
rect 622 278 626 282
rect 718 328 722 332
rect 734 358 738 362
rect 790 468 794 472
rect 758 458 762 462
rect 758 448 762 452
rect 782 448 786 452
rect 774 418 778 422
rect 774 408 778 412
rect 766 398 770 402
rect 814 468 818 472
rect 854 518 858 522
rect 838 508 842 512
rect 926 568 930 572
rect 966 668 970 672
rect 1002 903 1006 907
rect 1009 903 1013 907
rect 1070 948 1074 952
rect 1038 938 1042 942
rect 1054 938 1058 942
rect 1030 928 1034 932
rect 1062 878 1066 882
rect 1062 868 1066 872
rect 1038 848 1042 852
rect 1062 838 1066 842
rect 1022 788 1026 792
rect 990 748 994 752
rect 1014 728 1018 732
rect 982 708 986 712
rect 1002 703 1006 707
rect 1009 703 1013 707
rect 982 668 986 672
rect 990 648 994 652
rect 982 558 986 562
rect 910 548 914 552
rect 934 548 938 552
rect 886 538 890 542
rect 894 538 898 542
rect 950 538 954 542
rect 878 528 882 532
rect 934 528 938 532
rect 862 478 866 482
rect 878 478 882 482
rect 926 478 930 482
rect 886 468 890 472
rect 926 468 930 472
rect 814 438 818 442
rect 814 428 818 432
rect 798 388 802 392
rect 806 368 810 372
rect 750 348 754 352
rect 822 358 826 362
rect 974 548 978 552
rect 958 498 962 502
rect 974 498 978 502
rect 862 458 866 462
rect 918 458 922 462
rect 950 458 954 462
rect 854 448 858 452
rect 854 428 858 432
rect 870 428 874 432
rect 998 628 1002 632
rect 1102 938 1106 942
rect 1142 928 1146 932
rect 1094 918 1098 922
rect 1094 898 1098 902
rect 1158 918 1162 922
rect 1182 938 1186 942
rect 1198 938 1202 942
rect 1238 1068 1242 1072
rect 1406 1208 1410 1212
rect 1430 1188 1434 1192
rect 1478 1238 1482 1242
rect 1462 1168 1466 1172
rect 1454 1148 1458 1152
rect 1398 1138 1402 1142
rect 1406 1138 1410 1142
rect 1398 1128 1402 1132
rect 1414 1128 1418 1132
rect 1438 1128 1442 1132
rect 1302 1088 1306 1092
rect 1318 1088 1322 1092
rect 1302 1078 1306 1082
rect 1230 1058 1234 1062
rect 1246 1038 1250 1042
rect 1222 938 1226 942
rect 1222 928 1226 932
rect 1246 918 1250 922
rect 1174 908 1178 912
rect 1230 908 1234 912
rect 1286 898 1290 902
rect 1198 888 1202 892
rect 1182 878 1186 882
rect 1238 878 1242 882
rect 1246 878 1250 882
rect 1262 878 1266 882
rect 1078 868 1082 872
rect 1094 868 1098 872
rect 1110 868 1114 872
rect 1118 868 1122 872
rect 1158 868 1162 872
rect 1222 868 1226 872
rect 1174 858 1178 862
rect 1190 858 1194 862
rect 1142 838 1146 842
rect 1086 818 1090 822
rect 1078 798 1082 802
rect 1126 808 1130 812
rect 1070 788 1074 792
rect 1078 768 1082 772
rect 1086 758 1090 762
rect 1054 748 1058 752
rect 1062 748 1066 752
rect 1086 738 1090 742
rect 1046 728 1050 732
rect 1030 708 1034 712
rect 1054 718 1058 722
rect 1038 668 1042 672
rect 1046 648 1050 652
rect 1014 598 1018 602
rect 1006 578 1010 582
rect 1014 568 1018 572
rect 1014 548 1018 552
rect 1070 708 1074 712
rect 1062 658 1066 662
rect 1118 728 1122 732
rect 1110 708 1114 712
rect 1086 658 1090 662
rect 1118 678 1122 682
rect 1190 798 1194 802
rect 1230 858 1234 862
rect 1222 788 1226 792
rect 1206 768 1210 772
rect 1214 768 1218 772
rect 1142 758 1146 762
rect 1134 738 1138 742
rect 1190 738 1194 742
rect 1150 728 1154 732
rect 1238 818 1242 822
rect 1214 738 1218 742
rect 1230 738 1234 742
rect 1206 728 1210 732
rect 1198 718 1202 722
rect 1150 698 1154 702
rect 1166 698 1170 702
rect 1158 678 1162 682
rect 1174 678 1178 682
rect 1182 678 1186 682
rect 1126 668 1130 672
rect 1118 658 1122 662
rect 1126 648 1130 652
rect 1054 578 1058 582
rect 1118 608 1122 612
rect 1110 568 1114 572
rect 1086 558 1090 562
rect 1102 558 1106 562
rect 1062 548 1066 552
rect 1014 538 1018 542
rect 1038 538 1042 542
rect 1046 538 1050 542
rect 1030 528 1034 532
rect 1046 528 1050 532
rect 1158 658 1162 662
rect 1222 728 1226 732
rect 1254 868 1258 872
rect 1454 1098 1458 1102
rect 1470 1108 1474 1112
rect 1414 1068 1418 1072
rect 1422 1058 1426 1062
rect 1430 1058 1434 1062
rect 1462 1058 1466 1062
rect 1470 1058 1474 1062
rect 1398 1048 1402 1052
rect 1422 1048 1426 1052
rect 1399 958 1403 962
rect 1438 968 1442 972
rect 1478 958 1482 962
rect 1494 1198 1498 1202
rect 1438 948 1442 952
rect 1470 948 1474 952
rect 1486 948 1490 952
rect 1398 938 1402 942
rect 1454 928 1458 932
rect 1422 908 1426 912
rect 1302 888 1306 892
rect 1406 888 1410 892
rect 1310 878 1314 882
rect 1318 868 1322 872
rect 1262 858 1266 862
rect 1278 858 1282 862
rect 1286 828 1290 832
rect 1270 788 1274 792
rect 1286 768 1290 772
rect 1390 858 1394 862
rect 1398 858 1402 862
rect 1358 848 1362 852
rect 1374 848 1378 852
rect 1382 838 1386 842
rect 1358 798 1362 802
rect 1310 788 1314 792
rect 1318 788 1322 792
rect 1294 758 1298 762
rect 1302 758 1306 762
rect 1254 738 1258 742
rect 1302 738 1306 742
rect 1262 718 1266 722
rect 1302 708 1306 712
rect 1294 698 1298 702
rect 1286 688 1290 692
rect 1230 678 1234 682
rect 1238 678 1242 682
rect 1262 678 1266 682
rect 1206 668 1210 672
rect 1230 668 1234 672
rect 1254 668 1258 672
rect 1270 668 1274 672
rect 1190 658 1194 662
rect 1278 658 1282 662
rect 1166 648 1170 652
rect 1246 648 1250 652
rect 1278 648 1282 652
rect 1286 648 1290 652
rect 1254 638 1258 642
rect 1206 618 1210 622
rect 1230 618 1234 622
rect 1134 568 1138 572
rect 1150 568 1154 572
rect 1246 578 1250 582
rect 1190 558 1194 562
rect 1158 548 1162 552
rect 1206 548 1210 552
rect 1222 548 1226 552
rect 1230 548 1234 552
rect 1326 768 1330 772
rect 1342 768 1346 772
rect 1318 758 1322 762
rect 1366 778 1370 782
rect 1374 778 1378 782
rect 1374 758 1378 762
rect 1382 748 1386 752
rect 1390 748 1394 752
rect 1326 738 1330 742
rect 1358 738 1362 742
rect 1334 688 1338 692
rect 1318 668 1322 672
rect 1326 668 1330 672
rect 1366 668 1370 672
rect 1302 658 1306 662
rect 1350 658 1354 662
rect 1326 638 1330 642
rect 1326 578 1330 582
rect 1302 558 1306 562
rect 1358 618 1362 622
rect 1350 578 1354 582
rect 1294 548 1298 552
rect 1334 548 1338 552
rect 1374 638 1378 642
rect 1438 878 1442 882
rect 1446 878 1450 882
rect 1422 858 1426 862
rect 1478 848 1482 852
rect 1462 838 1466 842
rect 1502 838 1506 842
rect 1486 818 1490 822
rect 1454 758 1458 762
rect 1422 748 1426 752
rect 1430 738 1434 742
rect 1414 728 1418 732
rect 1398 698 1402 702
rect 1406 698 1410 702
rect 1438 698 1442 702
rect 1470 708 1474 712
rect 1462 688 1466 692
rect 1390 678 1394 682
rect 1382 558 1386 562
rect 1086 538 1090 542
rect 1262 538 1266 542
rect 1374 538 1378 542
rect 1094 528 1098 532
rect 1002 503 1006 507
rect 1009 503 1013 507
rect 1078 518 1082 522
rect 990 488 994 492
rect 1054 488 1058 492
rect 1038 478 1042 482
rect 990 468 994 472
rect 998 468 1002 472
rect 1014 468 1018 472
rect 974 458 978 462
rect 990 458 994 462
rect 1022 458 1026 462
rect 942 448 946 452
rect 958 448 962 452
rect 966 428 970 432
rect 886 418 890 422
rect 862 388 866 392
rect 918 388 922 392
rect 846 378 850 382
rect 838 368 842 372
rect 838 358 842 362
rect 814 348 818 352
rect 830 348 834 352
rect 846 348 850 352
rect 878 368 882 372
rect 870 358 874 362
rect 902 358 906 362
rect 798 338 802 342
rect 822 338 826 342
rect 830 338 834 342
rect 750 328 754 332
rect 742 318 746 322
rect 726 308 730 312
rect 750 308 754 312
rect 782 308 786 312
rect 694 288 698 292
rect 734 288 738 292
rect 678 278 682 282
rect 686 278 690 282
rect 590 258 594 262
rect 582 228 586 232
rect 614 268 618 272
rect 606 188 610 192
rect 702 278 706 282
rect 710 278 714 282
rect 670 258 674 262
rect 630 248 634 252
rect 686 248 690 252
rect 638 158 642 162
rect 598 148 602 152
rect 582 128 586 132
rect 582 98 586 102
rect 542 68 546 72
rect 558 68 562 72
rect 526 58 530 62
rect 542 58 546 62
rect 482 3 486 7
rect 489 3 493 7
rect 622 138 626 142
rect 654 238 658 242
rect 678 158 682 162
rect 774 288 778 292
rect 782 288 786 292
rect 790 288 794 292
rect 758 268 762 272
rect 814 298 818 302
rect 806 278 810 282
rect 942 378 946 382
rect 926 358 930 362
rect 910 348 914 352
rect 886 338 890 342
rect 918 338 922 342
rect 846 328 850 332
rect 886 328 890 332
rect 878 318 882 322
rect 870 298 874 302
rect 838 278 842 282
rect 862 278 866 282
rect 958 368 962 372
rect 1078 478 1082 482
rect 1062 468 1066 472
rect 1086 468 1090 472
rect 998 448 1002 452
rect 1014 448 1018 452
rect 1054 448 1058 452
rect 1086 448 1090 452
rect 1062 438 1066 442
rect 1046 428 1050 432
rect 1014 368 1018 372
rect 1086 398 1090 402
rect 1046 378 1050 382
rect 1078 378 1082 382
rect 1062 368 1066 372
rect 1046 358 1050 362
rect 1030 348 1034 352
rect 1046 348 1050 352
rect 1078 358 1082 362
rect 1086 358 1090 362
rect 1134 508 1138 512
rect 1118 488 1122 492
rect 1102 468 1106 472
rect 1102 378 1106 382
rect 1150 468 1154 472
rect 1190 528 1194 532
rect 1174 468 1178 472
rect 1158 448 1162 452
rect 1254 518 1258 522
rect 1294 518 1298 522
rect 1230 488 1234 492
rect 1214 468 1218 472
rect 1262 488 1266 492
rect 1270 488 1274 492
rect 1222 458 1226 462
rect 1366 518 1370 522
rect 1382 498 1386 502
rect 1342 478 1346 482
rect 1406 638 1410 642
rect 1422 628 1426 632
rect 1470 638 1474 642
rect 1454 618 1458 622
rect 1438 588 1442 592
rect 1454 548 1458 552
rect 1470 548 1474 552
rect 1494 548 1498 552
rect 1430 538 1434 542
rect 1462 538 1466 542
rect 1486 538 1490 542
rect 1430 528 1434 532
rect 1422 518 1426 522
rect 1414 508 1418 512
rect 1398 478 1402 482
rect 1318 468 1322 472
rect 1350 468 1354 472
rect 1366 468 1370 472
rect 1246 458 1250 462
rect 1278 458 1282 462
rect 1230 448 1234 452
rect 1174 428 1178 432
rect 1134 398 1138 402
rect 1126 388 1130 392
rect 1110 358 1114 362
rect 1230 438 1234 442
rect 1270 438 1274 442
rect 1238 408 1242 412
rect 1270 408 1274 412
rect 1214 398 1218 402
rect 1174 368 1178 372
rect 1094 348 1098 352
rect 1118 348 1122 352
rect 1150 348 1154 352
rect 1110 328 1114 332
rect 982 318 986 322
rect 1110 318 1114 322
rect 1002 303 1006 307
rect 1009 303 1013 307
rect 990 298 994 302
rect 1038 298 1042 302
rect 1126 298 1130 302
rect 1198 348 1202 352
rect 1182 328 1186 332
rect 1238 348 1242 352
rect 1206 308 1210 312
rect 1214 308 1218 312
rect 1286 378 1290 382
rect 1302 458 1306 462
rect 1366 448 1370 452
rect 1310 428 1314 432
rect 1398 448 1402 452
rect 1382 418 1386 422
rect 1294 328 1298 332
rect 1190 298 1194 302
rect 1222 298 1226 302
rect 1142 288 1146 292
rect 1150 288 1154 292
rect 1214 288 1218 292
rect 918 278 922 282
rect 958 278 962 282
rect 974 278 978 282
rect 1102 278 1106 282
rect 1158 278 1162 282
rect 894 268 898 272
rect 926 268 930 272
rect 710 258 714 262
rect 838 258 842 262
rect 942 268 946 272
rect 982 268 986 272
rect 1006 268 1010 272
rect 990 258 994 262
rect 758 248 762 252
rect 766 248 770 252
rect 742 188 746 192
rect 726 178 730 182
rect 750 168 754 172
rect 750 158 754 162
rect 662 148 666 152
rect 702 148 706 152
rect 670 138 674 142
rect 694 138 698 142
rect 726 138 730 142
rect 646 108 650 112
rect 638 88 642 92
rect 662 98 666 102
rect 606 78 610 82
rect 646 78 650 82
rect 678 128 682 132
rect 734 128 738 132
rect 694 118 698 122
rect 710 88 714 92
rect 854 248 858 252
rect 806 228 810 232
rect 806 218 810 222
rect 798 208 802 212
rect 774 198 778 202
rect 774 158 778 162
rect 854 158 858 162
rect 806 148 810 152
rect 766 138 770 142
rect 774 128 778 132
rect 702 78 706 82
rect 758 78 762 82
rect 686 68 690 72
rect 734 68 738 72
rect 590 18 594 22
rect 638 48 642 52
rect 662 48 666 52
rect 662 38 666 42
rect 598 8 602 12
rect 638 8 642 12
rect 710 58 714 62
rect 742 58 746 62
rect 726 48 730 52
rect 750 48 754 52
rect 686 8 690 12
rect 702 8 706 12
rect 782 88 786 92
rect 798 68 802 72
rect 790 58 794 62
rect 790 48 794 52
rect 862 128 866 132
rect 830 108 834 112
rect 854 108 858 112
rect 926 238 930 242
rect 886 218 890 222
rect 878 158 882 162
rect 942 228 946 232
rect 942 178 946 182
rect 982 178 986 182
rect 958 168 962 172
rect 902 148 906 152
rect 910 148 914 152
rect 918 128 922 132
rect 942 128 946 132
rect 894 108 898 112
rect 814 88 818 92
rect 822 88 826 92
rect 862 88 866 92
rect 910 78 914 82
rect 966 88 970 92
rect 1030 266 1034 270
rect 1054 268 1058 272
rect 1078 268 1082 272
rect 1118 268 1122 272
rect 1158 268 1162 272
rect 1070 248 1074 252
rect 1046 238 1050 242
rect 1070 228 1074 232
rect 1038 218 1042 222
rect 1038 198 1042 202
rect 990 138 994 142
rect 846 68 850 72
rect 862 68 866 72
rect 902 68 906 72
rect 918 68 922 72
rect 998 128 1002 132
rect 1002 103 1006 107
rect 1009 103 1013 107
rect 1006 78 1010 82
rect 1094 248 1098 252
rect 1166 258 1170 262
rect 1286 298 1290 302
rect 1270 278 1274 282
rect 1190 268 1194 272
rect 1238 268 1242 272
rect 1294 268 1298 272
rect 1414 428 1418 432
rect 1334 408 1338 412
rect 1358 408 1362 412
rect 1366 408 1370 412
rect 1406 408 1410 412
rect 1334 398 1338 402
rect 1382 358 1386 362
rect 1390 358 1394 362
rect 1342 348 1346 352
rect 1358 348 1362 352
rect 1374 348 1378 352
rect 1334 328 1338 332
rect 1318 318 1322 322
rect 1246 258 1250 262
rect 1262 258 1266 262
rect 1270 258 1274 262
rect 1134 238 1138 242
rect 1126 218 1130 222
rect 1118 208 1122 212
rect 1086 198 1090 202
rect 1062 168 1066 172
rect 1070 158 1074 162
rect 1102 158 1106 162
rect 1134 198 1138 202
rect 1142 178 1146 182
rect 1134 158 1138 162
rect 1054 138 1058 142
rect 1046 128 1050 132
rect 1150 168 1154 172
rect 1102 138 1106 142
rect 1094 128 1098 132
rect 1110 128 1114 132
rect 1118 128 1122 132
rect 1126 128 1130 132
rect 1078 118 1082 122
rect 1078 98 1082 102
rect 1102 108 1106 112
rect 1070 88 1074 92
rect 822 58 826 62
rect 926 58 930 62
rect 950 58 954 62
rect 1022 58 1026 62
rect 1038 58 1042 62
rect 1110 98 1114 102
rect 1198 248 1202 252
rect 1222 228 1226 232
rect 1262 218 1266 222
rect 1246 208 1250 212
rect 1230 198 1234 202
rect 1214 158 1218 162
rect 1150 98 1154 102
rect 1174 108 1178 112
rect 1302 258 1306 262
rect 1286 208 1290 212
rect 1270 188 1274 192
rect 1262 168 1266 172
rect 1286 168 1290 172
rect 1334 258 1338 262
rect 1326 188 1330 192
rect 1334 188 1338 192
rect 1382 328 1386 332
rect 1406 348 1410 352
rect 1406 338 1410 342
rect 1486 518 1490 522
rect 1478 498 1482 502
rect 1502 508 1506 512
rect 1494 498 1498 502
rect 1502 488 1506 492
rect 1478 478 1482 482
rect 1454 458 1458 462
rect 1438 368 1442 372
rect 1486 368 1490 372
rect 1430 348 1434 352
rect 1422 338 1426 342
rect 1478 338 1482 342
rect 1438 328 1442 332
rect 1398 288 1402 292
rect 1454 318 1458 322
rect 1366 268 1370 272
rect 1422 268 1426 272
rect 1390 258 1394 262
rect 1414 258 1418 262
rect 1342 178 1346 182
rect 1406 178 1410 182
rect 1358 168 1362 172
rect 1302 158 1306 162
rect 1366 158 1370 162
rect 1390 158 1394 162
rect 1206 118 1210 122
rect 1142 88 1146 92
rect 1166 88 1170 92
rect 1126 78 1130 82
rect 1078 58 1082 62
rect 1110 58 1114 62
rect 1366 138 1370 142
rect 1286 128 1290 132
rect 1342 128 1346 132
rect 1358 128 1362 132
rect 1310 118 1314 122
rect 1374 118 1378 122
rect 1294 88 1298 92
rect 1342 88 1346 92
rect 1222 78 1226 82
rect 1238 78 1242 82
rect 1246 78 1250 82
rect 1398 118 1402 122
rect 1454 268 1458 272
rect 1486 318 1490 322
rect 1486 278 1490 282
rect 1438 258 1442 262
rect 1502 258 1506 262
rect 1462 248 1466 252
rect 1430 228 1434 232
rect 1478 158 1482 162
rect 1494 148 1498 152
rect 1422 128 1426 132
rect 1414 108 1418 112
rect 1382 88 1386 92
rect 1430 108 1434 112
rect 1438 78 1442 82
rect 1462 78 1466 82
rect 1150 68 1154 72
rect 1182 68 1186 72
rect 1198 68 1202 72
rect 1238 68 1242 72
rect 1286 68 1290 72
rect 1366 68 1370 72
rect 1454 68 1458 72
rect 1486 68 1490 72
rect 1206 58 1210 62
rect 862 48 866 52
rect 886 48 890 52
rect 1022 48 1026 52
rect 1190 48 1194 52
rect 1206 48 1210 52
rect 1294 58 1298 62
rect 1318 58 1322 62
rect 1246 38 1250 42
rect 1374 58 1378 62
rect 1422 58 1426 62
rect 1462 58 1466 62
rect 1310 48 1314 52
rect 1334 48 1338 52
rect 1398 48 1402 52
rect 1254 18 1258 22
rect 1262 18 1266 22
<< metal3 >>
rect 1534 1321 1538 1322
rect 1522 1318 1538 1321
rect 1000 1303 1002 1307
rect 1006 1303 1009 1307
rect 1014 1303 1016 1307
rect 1534 1301 1538 1302
rect 1490 1298 1538 1301
rect 106 1288 462 1291
rect 138 1278 201 1281
rect 242 1278 270 1281
rect 402 1278 406 1281
rect 418 1278 566 1281
rect 626 1278 654 1281
rect 778 1278 790 1281
rect 914 1278 1102 1281
rect 1218 1278 1374 1281
rect 1534 1281 1538 1282
rect 1454 1278 1538 1281
rect 18 1268 38 1271
rect 70 1271 73 1278
rect 70 1268 142 1271
rect 154 1268 182 1271
rect 198 1271 201 1278
rect 198 1268 206 1271
rect 278 1271 281 1278
rect 1102 1272 1105 1278
rect 1454 1272 1457 1278
rect 210 1268 281 1271
rect 322 1268 414 1271
rect 458 1268 510 1271
rect 602 1268 638 1271
rect 650 1268 654 1271
rect 674 1268 686 1271
rect 738 1268 742 1271
rect 778 1268 846 1271
rect 6 1261 9 1268
rect 894 1262 897 1268
rect 6 1258 94 1261
rect 98 1258 118 1261
rect 162 1258 206 1261
rect 210 1258 305 1261
rect 314 1258 358 1261
rect 362 1258 398 1261
rect 402 1258 422 1261
rect 458 1258 502 1261
rect 618 1258 654 1261
rect 658 1258 718 1261
rect 722 1258 758 1261
rect 762 1258 806 1261
rect 954 1258 1030 1261
rect 1034 1258 1222 1261
rect 1534 1261 1538 1262
rect 1434 1258 1538 1261
rect 90 1248 94 1251
rect 126 1248 134 1251
rect 138 1248 174 1251
rect 242 1248 262 1251
rect 302 1251 305 1258
rect 302 1248 382 1251
rect 386 1248 550 1251
rect 562 1248 734 1251
rect 738 1248 814 1251
rect 818 1248 870 1251
rect 1034 1248 1438 1251
rect 1478 1242 1481 1248
rect 26 1238 38 1241
rect 42 1238 94 1241
rect 130 1238 230 1241
rect 258 1238 366 1241
rect 386 1238 406 1241
rect 418 1238 422 1241
rect 482 1238 510 1241
rect 514 1238 726 1241
rect 1534 1238 1538 1242
rect 702 1232 705 1238
rect 178 1228 270 1231
rect 298 1228 358 1231
rect 362 1228 446 1231
rect 450 1228 598 1231
rect 1406 1231 1409 1238
rect 1534 1231 1537 1238
rect 1406 1228 1537 1231
rect 194 1218 326 1221
rect 1002 1218 1414 1221
rect 34 1208 62 1211
rect 66 1208 382 1211
rect 554 1208 1126 1211
rect 1138 1208 1182 1211
rect 1186 1208 1406 1211
rect 480 1203 482 1207
rect 486 1203 489 1207
rect 494 1203 496 1207
rect 554 1198 598 1201
rect 650 1198 790 1201
rect 1170 1198 1278 1201
rect 1494 1192 1497 1198
rect 202 1188 558 1191
rect 590 1188 678 1191
rect 746 1188 1054 1191
rect 1074 1188 1086 1191
rect 590 1182 593 1188
rect 74 1178 238 1181
rect 346 1178 390 1181
rect 394 1178 422 1181
rect 426 1178 590 1181
rect 818 1178 1206 1181
rect 1430 1181 1433 1188
rect 1430 1178 1537 1181
rect 26 1168 38 1171
rect 42 1168 46 1171
rect 122 1168 150 1171
rect 270 1171 273 1178
rect 170 1168 257 1171
rect 270 1168 366 1171
rect 370 1168 430 1171
rect 718 1171 721 1178
rect 1534 1172 1537 1178
rect 718 1168 742 1171
rect 1018 1168 1094 1171
rect 1534 1168 1538 1172
rect 254 1162 257 1168
rect 1462 1162 1465 1168
rect 66 1158 110 1161
rect 130 1158 142 1161
rect 210 1158 222 1161
rect 306 1158 334 1161
rect 634 1158 670 1161
rect 1090 1158 1110 1161
rect 1130 1158 1142 1161
rect 1146 1158 1198 1161
rect 1218 1158 1286 1161
rect 50 1148 70 1151
rect 74 1148 150 1151
rect 154 1148 238 1151
rect 338 1148 358 1151
rect 362 1148 422 1151
rect 618 1148 662 1151
rect 674 1148 678 1151
rect 706 1148 750 1151
rect 754 1148 774 1151
rect 1050 1148 1094 1151
rect 1130 1148 1166 1151
rect 1178 1148 1198 1151
rect 1534 1151 1538 1152
rect 1458 1148 1538 1151
rect 22 1142 25 1148
rect 1206 1142 1209 1148
rect 34 1138 166 1141
rect 214 1138 286 1141
rect 322 1138 406 1141
rect 586 1138 606 1141
rect 650 1138 678 1141
rect 682 1138 734 1141
rect 1050 1138 1070 1141
rect 1074 1138 1142 1141
rect 1146 1138 1198 1141
rect 1402 1138 1406 1141
rect 214 1132 217 1138
rect 26 1128 54 1131
rect 114 1128 174 1131
rect 242 1128 294 1131
rect 298 1128 342 1131
rect 370 1128 398 1131
rect 546 1128 558 1131
rect 630 1131 633 1138
rect 630 1128 638 1131
rect 666 1128 694 1131
rect 698 1128 838 1131
rect 986 1128 1022 1131
rect 1186 1128 1398 1131
rect 1418 1128 1438 1131
rect 194 1118 302 1121
rect 346 1118 430 1121
rect 458 1118 558 1121
rect 602 1118 710 1121
rect 714 1118 806 1121
rect 962 1118 998 1121
rect 210 1108 270 1111
rect 322 1108 350 1111
rect 354 1108 566 1111
rect 818 1108 870 1111
rect 898 1108 926 1111
rect 318 1101 321 1108
rect 1000 1103 1002 1107
rect 1006 1103 1009 1107
rect 1014 1103 1016 1107
rect 1470 1102 1473 1108
rect 234 1098 321 1101
rect 330 1098 918 1101
rect 1114 1098 1454 1101
rect 90 1088 110 1091
rect 114 1088 169 1091
rect 258 1088 406 1091
rect 522 1088 606 1091
rect 626 1088 665 1091
rect 770 1088 862 1091
rect 866 1088 1001 1091
rect 1106 1088 1110 1091
rect 1114 1088 1302 1091
rect 1306 1088 1318 1091
rect 166 1082 169 1088
rect 662 1082 665 1088
rect 998 1082 1001 1088
rect 58 1078 126 1081
rect 202 1078 254 1081
rect 290 1078 350 1081
rect 514 1078 550 1081
rect 554 1078 646 1081
rect 714 1078 734 1081
rect 738 1078 785 1081
rect 914 1078 966 1081
rect 1218 1078 1302 1081
rect 782 1072 785 1078
rect 42 1068 86 1071
rect 90 1068 142 1071
rect 146 1068 158 1071
rect 162 1068 166 1071
rect 250 1068 326 1071
rect 346 1068 390 1071
rect 394 1068 438 1071
rect 442 1068 462 1071
rect 474 1068 510 1071
rect 562 1068 582 1071
rect 698 1068 718 1071
rect 722 1068 734 1071
rect 882 1068 886 1071
rect 1242 1068 1414 1071
rect 42 1058 78 1061
rect 178 1058 206 1061
rect 378 1058 382 1061
rect 410 1058 422 1061
rect 426 1058 454 1061
rect 474 1058 478 1061
rect 538 1058 582 1061
rect 586 1058 601 1061
rect 678 1061 681 1068
rect 634 1058 681 1061
rect 706 1058 742 1061
rect 746 1058 758 1061
rect 826 1058 830 1061
rect 922 1058 934 1061
rect 954 1058 974 1061
rect 978 1058 1038 1061
rect 1042 1058 1230 1061
rect 1426 1058 1430 1061
rect 1466 1058 1470 1061
rect 10 1048 14 1051
rect 66 1048 86 1051
rect 154 1048 182 1051
rect 298 1048 318 1051
rect 350 1051 353 1058
rect 598 1052 601 1058
rect 350 1048 382 1051
rect 434 1048 454 1051
rect 634 1048 638 1051
rect 650 1048 654 1051
rect 694 1051 697 1058
rect 674 1048 697 1051
rect 730 1048 750 1051
rect 754 1048 830 1051
rect 1162 1048 1198 1051
rect 1402 1048 1422 1051
rect 22 1041 25 1048
rect 22 1038 198 1041
rect 218 1038 230 1041
rect 266 1038 310 1041
rect 314 1038 318 1041
rect 330 1038 406 1041
rect 426 1038 478 1041
rect 550 1041 553 1048
rect 482 1038 553 1041
rect 562 1038 590 1041
rect 594 1038 622 1041
rect 818 1038 854 1041
rect 858 1038 910 1041
rect 1154 1038 1246 1041
rect 226 1028 246 1031
rect 282 1028 302 1031
rect 306 1028 334 1031
rect 338 1028 462 1031
rect 522 1028 534 1031
rect 538 1028 694 1031
rect 882 1028 1222 1031
rect 22 1022 25 1028
rect 562 1018 654 1021
rect 802 1018 838 1021
rect 842 1018 878 1021
rect 1202 1018 1214 1021
rect 514 1008 590 1011
rect 994 1008 1062 1011
rect 480 1003 482 1007
rect 486 1003 489 1007
rect 494 1003 496 1007
rect 82 988 102 991
rect 458 988 518 991
rect 826 988 862 991
rect 874 988 974 991
rect 1098 988 1198 991
rect 266 978 286 981
rect 290 978 318 981
rect 322 978 382 981
rect 474 978 518 981
rect 778 978 894 981
rect 970 978 1054 981
rect 26 968 54 971
rect 58 968 62 971
rect 90 968 166 971
rect 170 968 190 971
rect 346 968 398 971
rect 406 971 409 978
rect 402 968 430 971
rect 466 968 510 971
rect 514 968 542 971
rect 658 968 710 971
rect 714 968 790 971
rect 874 968 950 971
rect 1430 968 1438 971
rect 1534 971 1538 972
rect 1442 968 1538 971
rect 98 958 158 961
rect 162 958 206 961
rect 234 958 238 961
rect 378 958 542 961
rect 682 958 694 961
rect 746 958 766 961
rect 770 958 870 961
rect 990 961 993 968
rect 970 958 993 961
rect 1398 958 1399 961
rect 1482 958 1513 961
rect 50 948 62 951
rect 298 948 318 951
rect 362 948 390 951
rect 394 948 526 951
rect 626 948 718 951
rect 762 948 766 951
rect 778 948 790 951
rect 810 948 814 951
rect 822 948 918 951
rect 994 948 1070 951
rect 1398 951 1401 958
rect 1398 948 1438 951
rect 1442 948 1470 951
rect 1510 951 1513 958
rect 1534 951 1538 952
rect 1510 948 1538 951
rect 10 938 30 941
rect 126 938 222 941
rect 350 941 353 948
rect 250 938 353 941
rect 370 938 374 941
rect 394 938 406 941
rect 426 938 534 941
rect 538 938 550 941
rect 602 938 641 941
rect 650 938 670 941
rect 730 938 734 941
rect 778 938 782 941
rect 822 941 825 948
rect 1182 942 1185 948
rect 1486 942 1489 948
rect 786 938 825 941
rect 930 938 966 941
rect 1034 938 1038 941
rect 1058 938 1102 941
rect 1194 938 1198 941
rect 1226 938 1398 941
rect 126 932 129 938
rect 638 932 641 938
rect 1142 932 1145 938
rect 26 928 86 931
rect 90 928 118 931
rect 274 928 302 931
rect 306 928 502 931
rect 730 928 750 931
rect 754 928 830 931
rect 938 928 942 931
rect 946 928 990 931
rect 1034 928 1038 931
rect 1226 928 1454 931
rect 42 918 46 921
rect 254 921 257 928
rect 106 918 257 921
rect 338 918 438 921
rect 442 918 454 921
rect 530 918 550 921
rect 610 918 646 921
rect 714 918 766 921
rect 810 918 838 921
rect 850 918 910 921
rect 986 918 1094 921
rect 1162 918 1246 921
rect 162 908 254 911
rect 642 908 654 911
rect 698 908 718 911
rect 1178 908 1230 911
rect 1234 908 1422 911
rect 142 902 145 908
rect 1000 903 1002 907
rect 1006 903 1009 907
rect 1014 903 1016 907
rect 818 898 886 901
rect 890 898 945 901
rect 1098 898 1134 901
rect 1138 898 1286 901
rect 18 888 70 891
rect 162 888 214 891
rect 378 888 414 891
rect 450 888 542 891
rect 634 888 742 891
rect 882 888 934 891
rect 942 891 945 898
rect 942 888 1065 891
rect 82 878 102 881
rect 306 878 406 881
rect 410 878 566 881
rect 594 878 614 881
rect 618 878 638 881
rect 870 881 873 888
rect 1062 882 1065 888
rect 1306 888 1406 891
rect 870 878 942 881
rect 1198 881 1201 888
rect 1186 878 1201 881
rect 1242 878 1246 881
rect 1250 878 1262 881
rect 1266 878 1310 881
rect 1442 878 1446 881
rect 74 868 78 871
rect 90 868 126 871
rect 130 868 174 871
rect 258 868 270 871
rect 346 868 382 871
rect 402 868 406 871
rect 410 868 430 871
rect 490 868 534 871
rect 574 871 577 878
rect 862 872 865 878
rect 538 868 577 871
rect 610 868 742 871
rect 746 868 862 871
rect 914 868 1062 871
rect 1082 868 1094 871
rect 1122 868 1158 871
rect 1226 868 1238 871
rect 1258 868 1281 871
rect 1306 868 1318 871
rect 34 858 46 861
rect 50 858 94 861
rect 146 858 182 861
rect 282 858 326 861
rect 358 858 390 861
rect 426 858 470 861
rect 474 858 630 861
rect 762 858 814 861
rect 894 861 897 868
rect 818 858 897 861
rect 1110 861 1113 868
rect 1278 862 1281 868
rect 1110 858 1174 861
rect 1178 858 1190 861
rect 1194 858 1230 861
rect 1234 858 1262 861
rect 1358 858 1390 861
rect 1402 858 1422 861
rect 10 848 150 851
rect 202 848 254 851
rect 258 848 286 851
rect 298 848 318 851
rect 342 851 345 858
rect 322 848 345 851
rect 358 852 361 858
rect 390 852 393 858
rect 418 848 438 851
rect 442 848 446 851
rect 458 848 478 851
rect 482 848 526 851
rect 638 851 641 858
rect 1038 852 1041 858
rect 1358 852 1361 858
rect 570 848 641 851
rect 666 848 870 851
rect 1378 848 1465 851
rect 1534 851 1538 852
rect 1482 848 1538 851
rect 90 838 190 841
rect 194 838 329 841
rect 362 838 398 841
rect 534 841 537 848
rect 1462 842 1465 848
rect 522 838 537 841
rect 562 838 574 841
rect 602 838 646 841
rect 674 838 686 841
rect 858 838 1062 841
rect 1146 838 1358 841
rect 1362 838 1382 841
rect 1466 838 1502 841
rect 326 832 329 838
rect 854 832 857 838
rect 466 828 590 831
rect 594 828 614 831
rect 618 828 622 831
rect 634 828 854 831
rect 874 828 910 831
rect 914 828 934 831
rect 1290 828 1390 831
rect 98 818 126 821
rect 130 818 166 821
rect 170 818 174 821
rect 330 818 406 821
rect 410 818 566 821
rect 570 818 734 821
rect 738 818 766 821
rect 818 818 838 821
rect 882 818 958 821
rect 970 818 1086 821
rect 1242 818 1486 821
rect 538 808 550 811
rect 570 808 606 811
rect 738 808 758 811
rect 882 808 1126 811
rect 174 802 177 808
rect 480 803 482 807
rect 486 803 489 807
rect 494 803 496 807
rect 774 802 777 808
rect 514 798 558 801
rect 634 798 726 801
rect 730 798 750 801
rect 818 798 1078 801
rect 1082 798 1102 801
rect 1194 798 1358 801
rect 42 788 54 791
rect 82 788 142 791
rect 274 788 598 791
rect 722 788 734 791
rect 822 788 1022 791
rect 1074 788 1222 791
rect 1226 788 1270 791
rect 1274 788 1310 791
rect 1314 788 1318 791
rect 822 782 825 788
rect 458 778 494 781
rect 498 778 529 781
rect 526 772 529 778
rect 618 778 742 781
rect 746 778 806 781
rect 898 778 942 781
rect 1286 778 1366 781
rect 362 768 398 771
rect 434 768 502 771
rect 558 771 561 778
rect 1286 772 1289 778
rect 558 768 582 771
rect 690 768 758 771
rect 762 768 878 771
rect 890 768 918 771
rect 922 768 926 771
rect 962 768 1078 771
rect 1082 768 1206 771
rect 1374 771 1377 778
rect 1346 768 1377 771
rect 42 758 62 761
rect 106 758 126 761
rect 198 761 201 768
rect 178 758 201 761
rect 258 758 270 761
rect 334 761 337 768
rect 278 758 337 761
rect 378 758 406 761
rect 410 758 582 761
rect 586 758 782 761
rect 786 758 822 761
rect 850 758 854 761
rect 858 758 942 761
rect 954 758 974 761
rect 978 758 982 761
rect 1214 761 1217 768
rect 1146 758 1294 761
rect 1306 758 1318 761
rect 1326 761 1329 768
rect 1326 758 1366 761
rect 1370 758 1374 761
rect 66 748 70 751
rect 74 748 94 751
rect 210 748 230 751
rect 278 751 281 758
rect 990 752 993 758
rect 274 748 281 751
rect 314 748 358 751
rect 442 748 470 751
rect 506 748 542 751
rect 570 748 574 751
rect 626 748 662 751
rect 666 748 718 751
rect 754 748 806 751
rect 834 748 974 751
rect 1050 748 1054 751
rect 1086 751 1089 758
rect 1390 752 1393 758
rect 1066 748 1382 751
rect 1454 751 1457 758
rect 1426 748 1457 751
rect 82 738 134 741
rect 138 738 150 741
rect 194 738 225 741
rect 242 738 294 741
rect 338 738 390 741
rect 402 738 430 741
rect 434 738 454 741
rect 610 738 614 741
rect 730 738 902 741
rect 906 738 1086 741
rect 1130 738 1134 741
rect 1138 738 1190 741
rect 1218 738 1230 741
rect 1234 738 1254 741
rect 1306 738 1326 741
rect 1362 738 1430 741
rect 118 732 121 738
rect 182 732 185 738
rect 222 732 225 738
rect 526 732 529 738
rect 90 728 94 731
rect 170 728 174 731
rect 258 728 270 731
rect 346 728 422 731
rect 426 728 438 731
rect 594 728 814 731
rect 842 728 846 731
rect 946 728 1006 731
rect 1018 728 1046 731
rect 1122 728 1150 731
rect 1210 728 1222 731
rect 454 722 457 728
rect 218 718 254 721
rect 258 718 350 721
rect 370 718 446 721
rect 610 718 686 721
rect 698 718 702 721
rect 722 718 798 721
rect 802 718 830 721
rect 834 718 862 721
rect 918 721 921 728
rect 1414 722 1417 728
rect 918 718 950 721
rect 962 718 1046 721
rect 1058 718 1198 721
rect 1202 718 1262 721
rect 154 708 262 711
rect 394 708 398 711
rect 554 708 574 711
rect 658 708 774 711
rect 874 708 982 711
rect 1034 708 1054 711
rect 1074 708 1110 711
rect 1114 708 1302 711
rect 1306 708 1470 711
rect 1000 703 1002 707
rect 1006 703 1009 707
rect 1014 703 1016 707
rect 282 698 342 701
rect 354 698 366 701
rect 386 698 993 701
rect 1146 698 1150 701
rect 1170 698 1254 701
rect 1298 698 1398 701
rect 1410 698 1438 701
rect 10 688 49 691
rect 210 688 222 691
rect 226 688 302 691
rect 306 688 310 691
rect 314 688 358 691
rect 402 688 457 691
rect 562 688 614 691
rect 666 688 678 691
rect 690 688 750 691
rect 754 688 814 691
rect 826 688 854 691
rect 990 691 993 698
rect 990 688 1286 691
rect 1338 688 1462 691
rect 46 682 49 688
rect 454 682 457 688
rect 218 678 246 681
rect 250 678 286 681
rect 290 678 382 681
rect 586 678 630 681
rect 650 678 694 681
rect 706 678 710 681
rect 770 678 894 681
rect 898 678 942 681
rect 982 678 1118 681
rect 1162 678 1174 681
rect 1186 678 1230 681
rect 1242 678 1262 681
rect 1318 678 1390 681
rect -26 671 -22 672
rect -26 668 6 671
rect 90 668 110 671
rect 314 668 334 671
rect 354 668 366 671
rect 394 668 470 671
rect 550 671 553 678
rect 982 672 985 678
rect 1318 672 1321 678
rect 550 668 566 671
rect 626 668 670 671
rect 738 668 790 671
rect 846 668 942 671
rect 1042 668 1046 671
rect 1130 668 1206 671
rect 1258 668 1270 671
rect 1330 668 1366 671
rect 58 658 94 661
rect 146 658 158 661
rect 202 658 238 661
rect 642 658 742 661
rect 846 661 849 668
rect 786 658 849 661
rect 858 658 862 661
rect 882 658 902 661
rect 966 661 969 668
rect 1230 662 1233 668
rect 914 658 969 661
rect 1066 658 1086 661
rect 1122 658 1158 661
rect 1162 658 1190 661
rect 1282 658 1302 661
rect 1306 658 1350 661
rect 270 652 273 658
rect 10 648 22 651
rect 26 648 62 651
rect 90 648 102 651
rect 122 648 174 651
rect 290 648 326 651
rect 330 648 350 651
rect 402 648 526 651
rect 602 648 662 651
rect 666 648 702 651
rect 890 648 990 651
rect 1050 648 1126 651
rect 1170 648 1182 651
rect 1250 648 1278 651
rect 1282 648 1286 651
rect 1374 648 1409 651
rect 158 642 161 648
rect 286 642 289 648
rect 90 638 142 641
rect 170 638 190 641
rect 370 638 534 641
rect 538 638 598 641
rect 610 638 686 641
rect 702 641 705 648
rect 1374 642 1377 648
rect 1406 642 1409 648
rect 702 638 814 641
rect 818 638 878 641
rect 906 638 1014 641
rect 1082 638 1254 641
rect 1330 638 1334 641
rect 1442 638 1470 641
rect 82 628 262 631
rect 426 628 558 631
rect 642 628 726 631
rect 770 628 926 631
rect 1002 628 1422 631
rect 450 618 766 621
rect 802 618 822 621
rect 926 618 934 621
rect 938 618 1118 621
rect 1122 618 1206 621
rect 1234 618 1326 621
rect 1362 618 1454 621
rect 146 608 214 611
rect 554 608 606 611
rect 610 608 745 611
rect 754 608 1118 611
rect 480 603 482 607
rect 486 603 489 607
rect 494 603 496 607
rect 162 598 350 601
rect 562 598 622 601
rect 742 601 745 608
rect 742 598 814 601
rect 818 598 846 601
rect 850 598 910 601
rect 1018 598 1246 601
rect 458 588 486 591
rect 506 588 582 591
rect 986 588 1438 591
rect 246 581 249 588
rect 202 578 249 581
rect 546 578 630 581
rect 634 578 718 581
rect 810 578 894 581
rect 898 578 1006 581
rect 1058 578 1246 581
rect 1250 578 1326 581
rect 54 571 57 578
rect 50 568 57 571
rect 106 568 110 571
rect 234 568 254 571
rect 330 568 366 571
rect 378 568 694 571
rect 790 571 793 578
rect 790 568 926 571
rect 1050 568 1110 571
rect 1154 568 1262 571
rect 1350 571 1353 578
rect 1302 568 1353 571
rect 154 558 174 561
rect 194 558 318 561
rect 338 558 534 561
rect 538 558 598 561
rect 602 558 614 561
rect 674 558 750 561
rect 762 558 766 561
rect 818 558 870 561
rect 1014 561 1017 568
rect 1134 562 1137 568
rect 1302 562 1305 568
rect 986 558 1017 561
rect 1066 558 1086 561
rect 1106 558 1110 561
rect 1194 558 1225 561
rect 1222 552 1225 558
rect 1534 561 1538 562
rect 1386 558 1538 561
rect 1294 552 1297 558
rect 1334 552 1337 558
rect 42 548 102 551
rect 114 548 126 551
rect 226 548 262 551
rect 298 548 318 551
rect 322 548 358 551
rect 410 548 414 551
rect 426 548 454 551
rect 538 548 542 551
rect 610 548 646 551
rect 650 548 670 551
rect 722 548 726 551
rect 730 548 798 551
rect 914 548 934 551
rect 978 548 998 551
rect 1018 548 1062 551
rect 1066 548 1078 551
rect 1154 548 1158 551
rect 1210 548 1214 551
rect 1234 548 1238 551
rect 1458 548 1470 551
rect 1490 548 1494 551
rect 154 538 174 541
rect 242 538 246 541
rect 250 538 310 541
rect 390 541 393 548
rect 314 538 393 541
rect 434 538 542 541
rect 546 538 558 541
rect 674 538 686 541
rect 714 538 798 541
rect 890 538 894 541
rect 954 538 1014 541
rect 1050 538 1086 541
rect 1250 538 1262 541
rect 1378 538 1430 541
rect 606 532 609 538
rect 290 528 342 531
rect 346 528 465 531
rect 514 528 526 531
rect 530 528 534 531
rect 626 528 766 531
rect 770 528 830 531
rect 882 528 918 531
rect 922 528 934 531
rect 1026 528 1030 531
rect 1038 531 1041 538
rect 1462 532 1465 538
rect 1038 528 1046 531
rect 1082 528 1094 531
rect 1098 528 1190 531
rect 1254 528 1430 531
rect 1486 531 1489 538
rect 1474 528 1489 531
rect 462 522 465 528
rect 1254 522 1257 528
rect 10 518 158 521
rect 178 518 278 521
rect 298 518 326 521
rect 330 518 374 521
rect 522 518 550 521
rect 770 518 774 521
rect 826 518 854 521
rect 1074 518 1078 521
rect 1266 518 1294 521
rect 1298 518 1366 521
rect 1470 521 1473 528
rect 1426 518 1473 521
rect 1490 518 1494 521
rect 138 508 254 511
rect 442 508 518 511
rect 522 508 590 511
rect 698 508 702 511
rect 722 508 790 511
rect 842 508 982 511
rect 1058 508 1134 511
rect 1194 508 1414 511
rect 1498 508 1502 511
rect 1000 503 1002 507
rect 1006 503 1009 507
rect 1014 503 1016 507
rect 170 498 238 501
rect 474 498 542 501
rect 554 498 614 501
rect 634 498 838 501
rect 962 498 974 501
rect 1250 498 1382 501
rect 1482 498 1494 501
rect 74 488 94 491
rect 98 488 182 491
rect 186 488 678 491
rect 698 488 774 491
rect 826 488 974 491
rect 994 488 1054 491
rect 1234 488 1262 491
rect 1274 488 1414 491
rect 1482 488 1502 491
rect 1118 482 1121 488
rect 1262 482 1265 488
rect 82 478 110 481
rect 114 478 190 481
rect 274 478 358 481
rect 386 478 406 481
rect 410 478 438 481
rect 442 478 462 481
rect 498 478 502 481
rect 514 478 654 481
rect 658 478 694 481
rect 714 478 726 481
rect 754 478 862 481
rect 882 478 910 481
rect 930 478 1030 481
rect 1034 478 1038 481
rect 1046 478 1078 481
rect 1290 478 1342 481
rect 1402 478 1478 481
rect 1482 478 1494 481
rect 22 471 25 478
rect 22 468 38 471
rect 146 468 166 471
rect 314 468 438 471
rect 450 468 486 471
rect 546 468 582 471
rect 594 468 614 471
rect 618 468 638 471
rect 698 468 710 471
rect 802 468 814 471
rect 890 468 894 471
rect 930 468 990 471
rect 1002 468 1006 471
rect 1046 471 1049 478
rect 1018 468 1049 471
rect 1058 468 1062 471
rect 1090 468 1102 471
rect 1154 468 1174 471
rect 1218 468 1318 471
rect 1346 468 1350 471
rect 1354 468 1358 471
rect 86 462 89 468
rect 398 462 401 468
rect 534 462 537 468
rect 790 462 793 468
rect 1366 462 1369 468
rect 58 458 70 461
rect 178 458 190 461
rect 306 458 382 461
rect 386 458 390 461
rect 458 458 462 461
rect 482 458 510 461
rect 562 458 574 461
rect 626 458 670 461
rect 762 458 766 461
rect 810 458 862 461
rect 922 458 950 461
rect 978 458 990 461
rect 994 458 1022 461
rect 1026 458 1161 461
rect 1226 458 1246 461
rect 1282 458 1286 461
rect 1370 458 1454 461
rect 286 452 289 458
rect 1158 452 1161 458
rect 34 448 62 451
rect 66 448 145 451
rect 346 448 406 451
rect 466 448 518 451
rect 530 448 558 451
rect 658 448 662 451
rect 762 448 782 451
rect 858 448 942 451
rect 946 448 958 451
rect 1002 448 1014 451
rect 1058 448 1078 451
rect 1082 448 1086 451
rect 1302 451 1305 458
rect 1234 448 1305 451
rect 1370 448 1398 451
rect 142 442 145 448
rect 106 438 110 441
rect 282 438 310 441
rect 426 438 502 441
rect 518 441 521 448
rect 518 438 614 441
rect 690 438 718 441
rect 818 438 1062 441
rect 1066 438 1230 441
rect 1274 438 1294 441
rect 122 428 142 431
rect 346 428 526 431
rect 554 428 814 431
rect 858 428 870 431
rect 970 428 1046 431
rect 1178 428 1310 431
rect 1314 428 1414 431
rect 90 418 206 421
rect 418 418 758 421
rect 762 418 774 421
rect 778 418 886 421
rect 890 418 1382 421
rect 506 408 582 411
rect 586 408 622 411
rect 626 408 774 411
rect 1078 408 1238 411
rect 1258 408 1270 411
rect 1274 408 1334 411
rect 1338 408 1358 411
rect 1370 408 1406 411
rect 480 403 482 407
rect 486 403 489 407
rect 494 403 496 407
rect 522 398 598 401
rect 618 398 694 401
rect 706 398 726 401
rect 1078 401 1081 408
rect 770 398 1081 401
rect 1090 398 1134 401
rect 1162 398 1214 401
rect 1330 398 1334 401
rect 194 388 278 391
rect 398 388 550 391
rect 562 388 718 391
rect 722 388 798 391
rect 802 388 862 391
rect 866 388 918 391
rect 922 388 1126 391
rect 1202 388 1289 391
rect 398 382 401 388
rect 1286 382 1289 388
rect 154 378 214 381
rect 574 378 590 381
rect 610 378 846 381
rect 946 378 1046 381
rect 1050 378 1070 381
rect 1082 378 1102 381
rect 574 372 577 378
rect 186 368 206 371
rect 354 368 414 371
rect 602 368 806 371
rect 810 368 838 371
rect 882 368 958 371
rect 1018 368 1062 371
rect 1066 368 1174 371
rect 1442 368 1486 371
rect 78 362 81 368
rect 126 361 129 368
rect 126 358 254 361
rect 330 358 382 361
rect 738 358 822 361
rect 842 358 870 361
rect 906 358 926 361
rect 1050 358 1078 361
rect 1090 358 1110 361
rect 1386 358 1390 361
rect 1394 358 1438 361
rect 86 352 89 358
rect 26 348 30 351
rect 50 348 70 351
rect 106 348 166 351
rect 218 348 230 351
rect 378 348 478 351
rect 482 348 646 351
rect 706 348 710 351
rect 738 348 750 351
rect 822 348 830 351
rect 842 348 846 351
rect 866 348 910 351
rect 914 348 1030 351
rect 1050 348 1094 351
rect 1122 348 1150 351
rect 1202 348 1238 351
rect 1346 348 1358 351
rect 1362 348 1374 351
rect 1410 348 1430 351
rect 814 342 817 348
rect 822 342 825 348
rect 42 338 57 341
rect 66 338 78 341
rect 102 338 150 341
rect 162 338 366 341
rect 426 338 430 341
rect 434 338 462 341
rect 530 338 550 341
rect 554 338 558 341
rect 698 338 798 341
rect 834 338 886 341
rect 890 338 918 341
rect 922 338 1262 341
rect 1410 338 1422 341
rect 1426 338 1478 341
rect 54 332 57 338
rect 102 332 105 338
rect 178 328 206 331
rect 330 328 366 331
rect 658 328 718 331
rect 838 328 846 331
rect 850 328 886 331
rect 1114 328 1118 331
rect 1290 328 1294 331
rect 1338 328 1382 331
rect 1442 328 1462 331
rect 742 322 745 328
rect 750 322 753 328
rect 74 318 134 321
rect 146 318 190 321
rect 306 318 358 321
rect 362 318 526 321
rect 530 318 566 321
rect 570 318 646 321
rect 650 318 726 321
rect 882 318 982 321
rect 1098 318 1110 321
rect 1182 321 1185 328
rect 1182 318 1318 321
rect 1458 318 1486 321
rect 50 308 78 311
rect 82 308 102 311
rect 706 308 726 311
rect 754 308 782 311
rect 786 308 846 311
rect 1098 308 1206 311
rect 1210 308 1214 311
rect 1000 303 1002 307
rect 1006 303 1009 307
rect 1014 303 1016 307
rect 242 298 286 301
rect 450 298 606 301
rect 610 298 622 301
rect 650 298 814 301
rect 818 298 870 301
rect 962 298 990 301
rect 1042 298 1126 301
rect 1194 298 1222 301
rect 1226 298 1286 301
rect 10 288 158 291
rect 290 288 302 291
rect 386 288 406 291
rect 410 288 454 291
rect 458 288 462 291
rect 570 288 574 291
rect 594 288 654 291
rect 658 288 694 291
rect 738 288 774 291
rect 794 288 854 291
rect 862 288 1094 291
rect 1154 288 1174 291
rect 1218 288 1254 291
rect 1266 288 1398 291
rect 326 282 329 288
rect 58 278 94 281
rect 102 278 206 281
rect 394 278 502 281
rect 626 278 678 281
rect 690 278 702 281
rect 782 281 785 288
rect 862 282 865 288
rect 714 278 769 281
rect 782 278 806 281
rect 810 278 838 281
rect 922 278 958 281
rect 978 278 1094 281
rect 1142 281 1145 288
rect 1106 278 1145 281
rect 1162 278 1270 281
rect 1534 281 1538 282
rect 1490 278 1538 281
rect -26 271 -22 272
rect 102 271 105 278
rect -26 268 105 271
rect 138 268 174 271
rect 218 268 270 271
rect 306 268 414 271
rect 418 268 470 271
rect 618 268 734 271
rect 766 271 769 278
rect 766 268 894 271
rect 898 268 910 271
rect 946 268 950 271
rect 978 268 982 271
rect 1010 270 1033 271
rect 1010 268 1030 270
rect 26 258 70 261
rect 74 258 86 261
rect 166 258 182 261
rect 186 258 198 261
rect 210 258 254 261
rect 258 258 334 261
rect 426 258 446 261
rect 450 258 462 261
rect 566 261 569 268
rect 758 262 761 268
rect 566 258 574 261
rect 674 258 710 261
rect 834 258 838 261
rect 926 261 929 268
rect 1058 268 1062 271
rect 1082 268 1086 271
rect 1122 268 1126 271
rect 1154 268 1158 271
rect 1170 268 1190 271
rect 1234 268 1238 271
rect 1258 268 1273 271
rect 1298 268 1366 271
rect 1426 268 1454 271
rect 1270 262 1273 268
rect 926 258 990 261
rect 994 258 1166 261
rect 1250 258 1262 261
rect 1274 258 1302 261
rect 1306 258 1334 261
rect 1394 258 1414 261
rect 1442 258 1502 261
rect 1534 261 1538 262
rect 1506 258 1538 261
rect 166 252 169 258
rect 42 248 78 251
rect 82 248 118 251
rect 226 248 246 251
rect 250 248 310 251
rect 342 248 433 251
rect 442 248 518 251
rect 590 251 593 258
rect 766 252 769 258
rect 562 248 630 251
rect 690 248 750 251
rect 754 248 758 251
rect 858 248 1070 251
rect 1074 248 1094 251
rect 1178 248 1198 251
rect 1226 248 1462 251
rect 342 242 345 248
rect 430 242 433 248
rect 90 238 102 241
rect 162 238 198 241
rect 202 238 254 241
rect 434 238 534 241
rect 538 238 542 241
rect 658 238 822 241
rect 930 238 934 241
rect 1050 238 1134 241
rect 274 228 278 231
rect 514 228 582 231
rect 810 228 942 231
rect 1074 228 1222 231
rect 1226 228 1390 231
rect 1394 228 1430 231
rect 354 218 374 221
rect 570 218 742 221
rect 746 218 806 221
rect 890 218 1038 221
rect 1130 218 1262 221
rect 802 208 1078 211
rect 1082 208 1118 211
rect 1122 208 1246 211
rect 1266 208 1286 211
rect 480 203 482 207
rect 486 203 489 207
rect 494 203 496 207
rect 330 198 430 201
rect 778 198 1038 201
rect 1042 198 1086 201
rect 1138 198 1230 201
rect 186 188 201 191
rect 482 188 606 191
rect 610 188 622 191
rect 1086 191 1089 198
rect 1334 192 1337 198
rect 1086 188 1270 191
rect 1274 188 1326 191
rect 198 182 201 188
rect 18 178 153 181
rect 250 178 310 181
rect 314 178 326 181
rect 742 181 745 188
rect 730 178 745 181
rect 946 178 958 181
rect 986 178 1142 181
rect 1146 178 1214 181
rect 1218 178 1342 181
rect 1346 178 1406 181
rect 150 172 153 178
rect 342 171 345 178
rect 170 168 345 171
rect 370 168 398 171
rect 450 168 534 171
rect 754 168 926 171
rect 962 168 1062 171
rect 1154 168 1262 171
rect 1282 168 1286 171
rect 1290 168 1358 171
rect 62 161 65 168
rect 62 158 102 161
rect 146 158 166 161
rect 186 158 214 161
rect 282 158 318 161
rect 370 158 406 161
rect 410 158 438 161
rect 458 158 486 161
rect 558 161 561 168
rect 490 158 561 161
rect 642 158 678 161
rect 754 158 766 161
rect 778 158 854 161
rect 882 158 1062 161
rect 1074 158 1086 161
rect 1106 158 1134 161
rect 1218 158 1222 161
rect 1298 158 1302 161
rect 1370 158 1390 161
rect 1482 158 1486 161
rect 22 151 25 158
rect 38 151 41 158
rect 22 148 41 151
rect 66 148 134 151
rect 138 148 230 151
rect 234 148 294 151
rect 350 151 353 158
rect 298 148 353 151
rect 418 148 478 151
rect 506 148 550 151
rect 554 148 598 151
rect 602 148 654 151
rect 666 148 702 151
rect 810 148 830 151
rect 914 148 1342 151
rect 1346 148 1494 151
rect 66 138 190 141
rect 250 138 262 141
rect 306 138 318 141
rect 386 138 406 141
rect 466 138 510 141
rect 602 138 622 141
rect 626 138 670 141
rect 674 138 694 141
rect 730 138 766 141
rect 902 141 905 148
rect 902 138 990 141
rect 994 138 1054 141
rect 1066 138 1102 141
rect 1114 138 1286 141
rect 1290 138 1366 141
rect 1110 132 1113 138
rect 50 128 118 131
rect 122 128 238 131
rect 242 128 278 131
rect 282 128 494 131
rect 522 128 582 131
rect 586 128 678 131
rect 682 128 702 131
rect 730 128 734 131
rect 738 128 774 131
rect 866 128 918 131
rect 946 128 998 131
rect 1002 128 1046 131
rect 1050 128 1094 131
rect 1130 128 1246 131
rect 1250 128 1286 131
rect 1310 128 1342 131
rect 1362 128 1422 131
rect 98 118 126 121
rect 194 118 238 121
rect 242 118 350 121
rect 458 118 462 121
rect 698 118 1078 121
rect 1118 121 1121 128
rect 1310 122 1313 128
rect 1090 118 1121 121
rect 1210 118 1238 121
rect 1378 118 1398 121
rect 178 108 358 111
rect 362 108 390 111
rect 538 108 646 111
rect 834 108 854 111
rect 858 108 894 111
rect 1106 108 1174 111
rect 1418 108 1430 111
rect 1000 103 1002 107
rect 1006 103 1009 107
rect 1014 103 1016 107
rect 106 98 230 101
rect 234 98 286 101
rect 290 98 302 101
rect 354 98 358 101
rect 370 98 582 101
rect 666 98 977 101
rect 1082 98 1110 101
rect 1114 98 1150 101
rect 58 88 118 91
rect 122 88 182 91
rect 186 88 334 91
rect 338 88 638 91
rect 714 88 718 91
rect 818 88 822 91
rect 826 88 862 91
rect 882 88 966 91
rect 974 91 977 98
rect 974 88 1070 91
rect 1074 88 1142 91
rect 1146 88 1166 91
rect 1298 88 1342 91
rect 1346 88 1382 91
rect 34 78 62 81
rect 426 78 518 81
rect 522 78 606 81
rect 610 78 646 81
rect 706 78 758 81
rect 782 81 785 88
rect 782 78 894 81
rect 914 78 1006 81
rect 1010 78 1126 81
rect 1242 78 1246 81
rect 1282 78 1438 81
rect 1442 78 1462 81
rect 278 71 281 78
rect 374 71 377 78
rect 1222 72 1225 78
rect 278 68 377 71
rect 418 68 454 71
rect 458 68 494 71
rect 546 68 558 71
rect 690 68 734 71
rect 746 68 798 71
rect 802 68 846 71
rect 866 68 902 71
rect 922 68 942 71
rect 950 68 1110 71
rect 1114 68 1150 71
rect 1186 68 1198 71
rect 1242 68 1286 71
rect 1322 68 1366 71
rect 1458 68 1486 71
rect 950 62 953 68
rect 162 58 374 61
rect 378 58 398 61
rect 490 58 526 61
rect 546 58 558 61
rect 714 58 734 61
rect 746 58 790 61
rect 794 58 822 61
rect 826 58 926 61
rect 1026 58 1038 61
rect 1082 58 1110 61
rect 1210 58 1214 61
rect 1298 58 1318 61
rect 1378 58 1422 61
rect 1426 58 1462 61
rect 266 48 310 51
rect 626 48 638 51
rect 642 48 662 51
rect 730 48 750 51
rect 794 48 801 51
rect 866 48 878 51
rect 890 48 1022 51
rect 1026 48 1190 51
rect 1194 48 1206 51
rect 1210 48 1302 51
rect 1314 48 1318 51
rect 1338 48 1398 51
rect 666 38 1246 41
rect 594 18 1254 21
rect 1258 18 1262 21
rect 274 8 278 11
rect 602 8 638 11
rect 690 8 702 11
rect 480 3 482 7
rect 486 3 489 7
rect 494 3 496 7
<< m4contact >>
rect 1002 1303 1006 1307
rect 1010 1303 1013 1307
rect 1013 1303 1014 1307
rect 398 1278 402 1282
rect 414 1278 418 1282
rect 1102 1278 1106 1282
rect 654 1268 658 1272
rect 734 1268 738 1272
rect 894 1268 898 1272
rect 870 1248 874 1252
rect 1478 1248 1482 1252
rect 406 1238 410 1242
rect 422 1238 426 1242
rect 326 1218 330 1222
rect 1126 1208 1130 1212
rect 482 1203 486 1207
rect 490 1203 493 1207
rect 493 1203 494 1207
rect 1494 1188 1498 1192
rect 238 1178 242 1182
rect 1206 1178 1210 1182
rect 46 1168 50 1172
rect 142 1158 146 1162
rect 1462 1158 1466 1162
rect 22 1148 26 1152
rect 1094 1148 1098 1152
rect 1126 1148 1130 1152
rect 1198 1148 1202 1152
rect 1206 1138 1210 1142
rect 22 1128 26 1132
rect 558 1118 562 1122
rect 894 1108 898 1112
rect 1002 1103 1006 1107
rect 1010 1103 1013 1107
rect 1013 1103 1014 1107
rect 326 1098 330 1102
rect 1470 1098 1474 1102
rect 1102 1088 1106 1092
rect 158 1068 162 1072
rect 326 1068 330 1072
rect 886 1068 890 1072
rect 382 1058 386 1062
rect 470 1058 474 1062
rect 934 1058 938 1062
rect 6 1048 10 1052
rect 630 1048 634 1052
rect 654 1048 658 1052
rect 310 1038 314 1042
rect 422 1038 426 1042
rect 558 1038 562 1042
rect 22 1028 26 1032
rect 1222 1028 1226 1032
rect 990 1008 994 1012
rect 482 1003 486 1007
rect 490 1003 493 1007
rect 493 1003 494 1007
rect 870 988 874 992
rect 62 968 66 972
rect 238 958 242 962
rect 526 948 530 952
rect 1182 948 1186 952
rect 374 938 378 942
rect 390 938 394 942
rect 550 938 554 942
rect 734 938 738 942
rect 774 938 778 942
rect 1030 938 1034 942
rect 1142 938 1146 942
rect 1190 938 1194 942
rect 1486 938 1490 942
rect 942 928 946 932
rect 1038 928 1042 932
rect 46 918 50 922
rect 526 918 530 922
rect 142 908 146 912
rect 158 908 162 912
rect 654 908 658 912
rect 1002 903 1006 907
rect 1010 903 1013 907
rect 1013 903 1014 907
rect 1134 898 1138 902
rect 566 878 570 882
rect 638 878 642 882
rect 78 868 82 872
rect 406 868 410 872
rect 862 868 866 872
rect 1238 868 1242 872
rect 1302 868 1306 872
rect 326 858 330 862
rect 1038 858 1042 862
rect 390 848 394 852
rect 414 848 418 852
rect 454 848 458 852
rect 566 848 570 852
rect 398 838 402 842
rect 1358 838 1362 842
rect 622 828 626 832
rect 854 828 858 832
rect 1390 828 1394 832
rect 174 818 178 822
rect 766 818 770 822
rect 814 818 818 822
rect 566 808 570 812
rect 774 808 778 812
rect 878 808 882 812
rect 482 803 486 807
rect 490 803 493 807
rect 493 803 494 807
rect 174 798 178 802
rect 1102 798 1106 802
rect 734 788 738 792
rect 806 778 810 782
rect 878 768 882 772
rect 926 768 930 772
rect 62 758 66 762
rect 942 758 946 762
rect 982 758 986 762
rect 990 758 994 762
rect 1366 758 1370 762
rect 1390 758 1394 762
rect 70 748 74 752
rect 310 748 314 752
rect 718 748 722 752
rect 1046 748 1050 752
rect 182 738 186 742
rect 238 738 242 742
rect 526 738 530 742
rect 614 738 618 742
rect 1126 738 1130 742
rect 174 728 178 732
rect 454 728 458 732
rect 590 728 594 732
rect 846 728 850 732
rect 1006 728 1010 732
rect 366 718 370 722
rect 702 718 706 722
rect 1046 718 1050 722
rect 1414 718 1418 722
rect 390 708 394 712
rect 550 708 554 712
rect 774 708 778 712
rect 1054 708 1058 712
rect 1002 703 1006 707
rect 1010 703 1013 707
rect 1013 703 1014 707
rect 1142 698 1146 702
rect 1254 698 1258 702
rect 6 688 10 692
rect 398 688 402 692
rect 686 688 690 692
rect 814 688 818 692
rect 854 688 858 692
rect 694 678 698 682
rect 766 678 770 682
rect 6 668 10 672
rect 350 668 354 672
rect 566 668 570 672
rect 1046 668 1050 672
rect 270 658 274 662
rect 862 658 866 662
rect 1230 658 1234 662
rect 286 648 290 652
rect 1182 648 1186 652
rect 166 638 170 642
rect 598 638 602 642
rect 606 638 610 642
rect 1014 638 1018 642
rect 1078 638 1082 642
rect 1334 638 1338 642
rect 1438 638 1442 642
rect 822 618 826 622
rect 1118 618 1122 622
rect 1326 618 1330 622
rect 550 608 554 612
rect 482 603 486 607
rect 490 603 493 607
rect 493 603 494 607
rect 558 598 562 602
rect 814 598 818 602
rect 1246 598 1250 602
rect 982 588 986 592
rect 542 578 546 582
rect 894 578 898 582
rect 110 568 114 572
rect 694 568 698 572
rect 1046 568 1050 572
rect 1262 568 1266 572
rect 534 558 538 562
rect 766 558 770 562
rect 1062 558 1066 562
rect 1110 558 1114 562
rect 1134 558 1138 562
rect 1294 558 1298 562
rect 1334 558 1338 562
rect 414 548 418 552
rect 542 548 546 552
rect 718 548 722 552
rect 998 548 1002 552
rect 1078 548 1082 552
rect 1150 548 1154 552
rect 1214 548 1218 552
rect 1238 548 1242 552
rect 1486 548 1490 552
rect 558 538 562 542
rect 606 538 610 542
rect 686 538 690 542
rect 798 538 802 542
rect 1246 538 1250 542
rect 622 528 626 532
rect 830 528 834 532
rect 918 528 922 532
rect 1022 528 1026 532
rect 1078 528 1082 532
rect 1462 528 1466 532
rect 1470 528 1474 532
rect 774 518 778 522
rect 822 518 826 522
rect 1070 518 1074 522
rect 1262 518 1266 522
rect 1494 518 1498 522
rect 694 508 698 512
rect 982 508 986 512
rect 1054 508 1058 512
rect 1190 508 1194 512
rect 1494 508 1498 512
rect 1002 503 1006 507
rect 1010 503 1013 507
rect 1013 503 1014 507
rect 838 498 842 502
rect 1246 498 1250 502
rect 974 488 978 492
rect 1414 488 1418 492
rect 1478 488 1482 492
rect 502 478 506 482
rect 710 478 714 482
rect 910 478 914 482
rect 1030 478 1034 482
rect 1118 478 1122 482
rect 1262 478 1266 482
rect 1286 478 1290 482
rect 1494 478 1498 482
rect 446 468 450 472
rect 534 468 538 472
rect 798 468 802 472
rect 894 468 898 472
rect 1006 468 1010 472
rect 1054 468 1058 472
rect 1342 468 1346 472
rect 1358 468 1362 472
rect 86 458 90 462
rect 286 458 290 462
rect 390 458 394 462
rect 454 458 458 462
rect 558 458 562 462
rect 766 458 770 462
rect 790 458 794 462
rect 806 458 810 462
rect 1286 458 1290 462
rect 1366 458 1370 462
rect 654 448 658 452
rect 1078 448 1082 452
rect 102 438 106 442
rect 502 438 506 442
rect 718 438 722 442
rect 1294 438 1298 442
rect 414 418 418 422
rect 758 418 762 422
rect 502 408 506 412
rect 1254 408 1258 412
rect 482 403 486 407
rect 490 403 493 407
rect 493 403 494 407
rect 694 398 698 402
rect 726 398 730 402
rect 1158 398 1162 402
rect 1326 398 1330 402
rect 550 388 554 392
rect 1198 388 1202 392
rect 590 378 594 382
rect 606 378 610 382
rect 1070 378 1074 382
rect 78 358 82 362
rect 86 358 90 362
rect 326 358 330 362
rect 1438 358 1442 362
rect 22 348 26 352
rect 102 348 106 352
rect 646 348 650 352
rect 702 348 706 352
rect 734 348 738 352
rect 838 348 842 352
rect 862 348 866 352
rect 366 338 370 342
rect 422 338 426 342
rect 550 338 554 342
rect 814 338 818 342
rect 1262 338 1266 342
rect 742 328 746 332
rect 1118 328 1122 332
rect 1286 328 1290 332
rect 1462 328 1466 332
rect 726 318 730 322
rect 750 318 754 322
rect 1094 318 1098 322
rect 78 308 82 312
rect 702 308 706 312
rect 846 308 850 312
rect 1094 308 1098 312
rect 1002 303 1006 307
rect 1010 303 1013 307
rect 1013 303 1014 307
rect 606 298 610 302
rect 958 298 962 302
rect 326 288 330 292
rect 462 288 466 292
rect 566 288 570 292
rect 854 288 858 292
rect 1094 288 1098 292
rect 1174 288 1178 292
rect 1254 288 1258 292
rect 1262 288 1266 292
rect 502 278 506 282
rect 1094 278 1098 282
rect 270 268 274 272
rect 414 268 418 272
rect 734 268 738 272
rect 910 268 914 272
rect 950 268 954 272
rect 974 268 978 272
rect 574 258 578 262
rect 758 258 762 262
rect 766 258 770 262
rect 830 258 834 262
rect 1062 268 1066 272
rect 1086 268 1090 272
rect 1126 268 1130 272
rect 1150 268 1154 272
rect 1166 268 1170 272
rect 1230 268 1234 272
rect 1254 268 1258 272
rect 310 248 314 252
rect 750 248 754 252
rect 1174 248 1178 252
rect 1222 248 1226 252
rect 542 238 546 242
rect 822 238 826 242
rect 934 238 938 242
rect 270 228 274 232
rect 1390 228 1394 232
rect 350 218 354 222
rect 742 218 746 222
rect 1078 208 1082 212
rect 1262 208 1266 212
rect 482 203 486 207
rect 490 203 493 207
rect 493 203 494 207
rect 1334 198 1338 202
rect 622 188 626 192
rect 958 178 962 182
rect 1214 178 1218 182
rect 926 168 930 172
rect 1262 168 1266 172
rect 1278 168 1282 172
rect 454 158 458 162
rect 766 158 770 162
rect 1062 158 1066 162
rect 1086 158 1090 162
rect 1222 158 1226 162
rect 1294 158 1298 162
rect 1486 158 1490 162
rect 654 148 658 152
rect 830 148 834 152
rect 1342 148 1346 152
rect 598 138 602 142
rect 1062 138 1066 142
rect 1110 138 1114 142
rect 1286 138 1290 142
rect 702 128 706 132
rect 726 128 730 132
rect 1246 128 1250 132
rect 350 118 354 122
rect 454 118 458 122
rect 1086 118 1090 122
rect 1238 118 1242 122
rect 1002 103 1006 107
rect 1010 103 1013 107
rect 1013 103 1014 107
rect 358 98 362 102
rect 366 98 370 102
rect 718 88 722 92
rect 878 88 882 92
rect 422 78 426 82
rect 894 78 898 82
rect 1278 78 1282 82
rect 742 68 746 72
rect 942 68 946 72
rect 1110 68 1114 72
rect 1222 68 1226 72
rect 1318 68 1322 72
rect 558 58 562 62
rect 734 58 738 62
rect 1214 58 1218 62
rect 622 48 626 52
rect 878 48 882 52
rect 1302 48 1306 52
rect 1318 48 1322 52
rect 278 8 282 12
rect 482 3 486 7
rect 490 3 493 7
rect 493 3 494 7
<< metal4 >>
rect 1000 1303 1002 1307
rect 1006 1303 1009 1307
rect 1014 1303 1016 1307
rect 402 1278 409 1281
rect 406 1242 409 1278
rect 414 1241 417 1278
rect 658 1268 662 1271
rect 738 1268 742 1271
rect 414 1238 422 1241
rect 22 1132 25 1148
rect 6 692 9 1048
rect 22 1032 25 1128
rect 46 922 49 1168
rect 62 762 65 968
rect 142 912 145 1158
rect 158 912 161 1068
rect 238 962 241 1178
rect 326 1102 329 1218
rect 480 1203 482 1207
rect 486 1203 489 1207
rect 494 1203 496 1207
rect 330 1068 334 1071
rect 378 1058 382 1061
rect 466 1058 470 1061
rect 558 1042 561 1118
rect 634 1048 641 1051
rect 314 1038 318 1041
rect 418 1038 422 1041
rect 480 1003 482 1007
rect 486 1003 489 1007
rect 494 1003 496 1007
rect 366 938 374 941
rect 70 868 78 871
rect 70 752 73 868
rect 326 852 329 858
rect 166 818 174 821
rect 10 668 14 671
rect 166 642 169 818
rect 174 732 177 798
rect 186 738 190 741
rect 234 738 238 741
rect 102 568 110 571
rect 86 362 89 458
rect 102 442 105 568
rect 26 348 30 351
rect 78 312 81 358
rect 98 348 102 351
rect 270 272 273 658
rect 286 462 289 648
rect 310 252 313 748
rect 366 722 369 938
rect 390 852 393 938
rect 526 922 529 948
rect 398 868 406 871
rect 390 712 393 848
rect 398 842 401 868
rect 410 848 414 851
rect 398 692 401 838
rect 454 732 457 848
rect 480 803 482 807
rect 486 803 489 807
rect 494 803 496 807
rect 526 742 529 918
rect 550 712 553 938
rect 638 882 641 1048
rect 654 912 657 1048
rect 870 992 873 1248
rect 894 1112 897 1268
rect 1000 1103 1002 1107
rect 1006 1103 1009 1107
rect 1014 1103 1016 1107
rect 882 1068 886 1071
rect 566 852 569 878
rect 566 672 569 808
rect 606 738 614 741
rect 346 668 350 671
rect 480 603 482 607
rect 486 603 489 607
rect 494 603 496 607
rect 394 458 398 461
rect 414 422 417 548
rect 506 478 510 481
rect 446 462 449 468
rect 326 292 329 358
rect 270 11 273 228
rect 350 122 353 218
rect 350 101 353 118
rect 366 102 369 338
rect 414 272 417 418
rect 350 98 358 101
rect 422 82 425 338
rect 454 162 457 458
rect 502 442 505 478
rect 534 472 537 558
rect 542 552 545 578
rect 480 403 482 407
rect 486 403 489 407
rect 494 403 496 407
rect 462 121 465 288
rect 502 282 505 408
rect 542 242 545 548
rect 550 392 553 608
rect 558 542 561 598
rect 558 462 561 538
rect 554 338 561 341
rect 480 203 482 207
rect 486 203 489 207
rect 494 203 496 207
rect 458 118 465 121
rect 558 62 561 338
rect 566 292 569 668
rect 590 382 593 728
rect 606 642 609 738
rect 578 258 582 261
rect 598 142 601 638
rect 606 382 609 538
rect 622 532 625 828
rect 734 792 737 938
rect 694 718 702 721
rect 686 542 689 688
rect 694 682 697 718
rect 694 572 697 678
rect 694 512 697 568
rect 718 552 721 748
rect 766 682 769 818
rect 774 812 777 938
rect 706 478 710 481
rect 606 302 609 378
rect 646 352 649 428
rect 622 52 625 188
rect 654 152 657 448
rect 694 402 697 468
rect 766 462 769 558
rect 774 522 777 708
rect 798 532 801 538
rect 706 348 710 351
rect 702 132 705 308
rect 718 92 721 438
rect 726 322 729 398
rect 726 132 729 318
rect 734 272 737 348
rect 742 222 745 328
rect 750 252 753 318
rect 758 262 761 418
rect 774 261 777 518
rect 794 468 798 471
rect 806 462 809 778
rect 814 692 817 818
rect 838 728 846 731
rect 814 672 817 688
rect 794 458 798 461
rect 814 342 817 598
rect 822 522 825 618
rect 770 258 777 261
rect 766 162 769 258
rect 822 242 825 518
rect 830 262 833 528
rect 838 502 841 728
rect 854 692 857 828
rect 862 662 865 868
rect 878 772 881 808
rect 918 768 926 771
rect 894 472 897 578
rect 918 532 921 768
rect 914 478 918 481
rect 842 348 849 351
rect 858 348 862 351
rect 846 312 849 348
rect 854 282 857 288
rect 914 268 918 271
rect 830 152 833 258
rect 934 242 937 1058
rect 942 762 945 928
rect 990 762 993 1008
rect 1000 903 1002 907
rect 1006 903 1009 907
rect 1014 903 1016 907
rect 982 592 985 758
rect 1006 732 1009 738
rect 1000 703 1002 707
rect 1006 703 1009 707
rect 1014 703 1016 707
rect 1018 638 1022 641
rect 974 492 977 558
rect 1002 548 1006 551
rect 1018 528 1022 531
rect 982 472 985 508
rect 1000 503 1002 507
rect 1006 503 1009 507
rect 1014 503 1016 507
rect 1030 482 1033 938
rect 1038 862 1041 928
rect 1046 722 1049 748
rect 1042 668 1046 671
rect 1046 572 1049 668
rect 1054 512 1057 708
rect 1074 638 1078 641
rect 1054 472 1057 478
rect 1006 462 1009 468
rect 1000 303 1002 307
rect 1006 303 1009 307
rect 1014 303 1016 307
rect 946 268 950 271
rect 958 182 961 298
rect 974 272 977 278
rect 1062 272 1065 558
rect 1078 532 1081 548
rect 1070 382 1073 518
rect 1082 448 1089 451
rect 1086 432 1089 448
rect 1094 322 1097 1148
rect 1102 1092 1105 1278
rect 1126 1152 1129 1208
rect 1102 561 1105 798
rect 1122 738 1126 741
rect 1102 558 1110 561
rect 1110 331 1113 558
rect 1118 482 1121 618
rect 1134 562 1137 898
rect 1142 702 1145 938
rect 1182 652 1185 948
rect 1110 328 1118 331
rect 1094 292 1097 308
rect 1150 282 1153 548
rect 1190 512 1193 938
rect 1078 268 1086 271
rect 1078 212 1081 268
rect 1094 192 1097 278
rect 1122 268 1126 271
rect 1158 271 1161 398
rect 1198 392 1201 1148
rect 1206 1142 1209 1178
rect 1210 548 1214 551
rect 1154 268 1161 271
rect 1166 272 1169 278
rect 1158 262 1161 268
rect 1174 252 1177 288
rect 1222 252 1225 1028
rect 1242 868 1246 871
rect 1298 868 1302 871
rect 1230 272 1233 658
rect 1238 532 1241 548
rect 1246 542 1249 598
rect 1246 502 1249 538
rect 1234 268 1241 271
rect 930 168 934 171
rect 1062 142 1065 158
rect 1086 122 1089 158
rect 1000 103 1002 107
rect 1006 103 1009 107
rect 1014 103 1016 107
rect 742 61 745 68
rect 738 58 745 61
rect 878 52 881 88
rect 898 78 902 81
rect 1110 72 1113 138
rect 942 52 945 68
rect 1214 62 1217 178
rect 1222 162 1225 168
rect 1222 72 1225 158
rect 1238 122 1241 268
rect 1246 132 1249 498
rect 1254 412 1257 698
rect 1326 638 1334 641
rect 1326 622 1329 638
rect 1262 522 1265 568
rect 1262 342 1265 478
rect 1286 472 1289 478
rect 1286 462 1289 468
rect 1294 442 1297 558
rect 1262 292 1265 338
rect 1254 272 1257 288
rect 1262 172 1265 208
rect 1274 168 1278 171
rect 1286 142 1289 328
rect 1294 162 1297 438
rect 1326 402 1329 618
rect 1334 552 1337 558
rect 1358 472 1361 838
rect 1390 762 1393 828
rect 1334 192 1337 198
rect 1298 158 1305 161
rect 1274 78 1278 81
rect 1302 52 1305 158
rect 1342 152 1345 468
rect 1366 462 1369 758
rect 1390 232 1393 758
rect 1414 492 1417 718
rect 1438 362 1441 638
rect 1462 532 1465 1158
rect 1470 532 1473 1098
rect 1462 332 1465 528
rect 1478 492 1481 1248
rect 1486 552 1489 938
rect 1486 162 1489 548
rect 1494 522 1497 1188
rect 1494 482 1497 508
rect 1318 52 1321 68
rect 1314 48 1318 51
rect 270 8 278 11
rect 480 3 482 7
rect 486 3 489 7
rect 494 3 496 7
<< m5contact >>
rect 1002 1303 1006 1307
rect 1009 1303 1010 1307
rect 1010 1303 1013 1307
rect 662 1268 666 1272
rect 742 1268 746 1272
rect 482 1203 486 1207
rect 489 1203 490 1207
rect 490 1203 493 1207
rect 334 1068 338 1072
rect 374 1058 378 1062
rect 462 1058 466 1062
rect 318 1038 322 1042
rect 414 1038 418 1042
rect 482 1003 486 1007
rect 489 1003 490 1007
rect 490 1003 493 1007
rect 326 848 330 852
rect 14 668 18 672
rect 190 738 194 742
rect 230 738 234 742
rect 30 348 34 352
rect 94 348 98 352
rect 406 848 410 852
rect 482 803 486 807
rect 489 803 490 807
rect 490 803 493 807
rect 1002 1103 1006 1107
rect 1009 1103 1010 1107
rect 1010 1103 1013 1107
rect 878 1068 882 1072
rect 342 668 346 672
rect 482 603 486 607
rect 489 603 490 607
rect 490 603 493 607
rect 398 458 402 462
rect 510 478 514 482
rect 446 458 450 462
rect 482 403 486 407
rect 489 403 490 407
rect 490 403 493 407
rect 482 203 486 207
rect 489 203 490 207
rect 490 203 493 207
rect 582 258 586 262
rect 702 478 706 482
rect 694 468 698 472
rect 646 428 650 432
rect 798 528 802 532
rect 710 348 714 352
rect 790 468 794 472
rect 814 668 818 672
rect 798 458 802 462
rect 918 478 922 482
rect 854 348 858 352
rect 854 278 858 282
rect 918 268 922 272
rect 1002 903 1006 907
rect 1009 903 1010 907
rect 1010 903 1013 907
rect 1006 738 1010 742
rect 1002 703 1006 707
rect 1009 703 1010 707
rect 1010 703 1013 707
rect 1022 638 1026 642
rect 974 558 978 562
rect 1006 548 1010 552
rect 1014 528 1018 532
rect 1002 503 1006 507
rect 1009 503 1010 507
rect 1010 503 1013 507
rect 1038 668 1042 672
rect 1070 638 1074 642
rect 1054 478 1058 482
rect 982 468 986 472
rect 1006 458 1010 462
rect 1002 303 1006 307
rect 1009 303 1010 307
rect 1010 303 1013 307
rect 942 268 946 272
rect 974 278 978 282
rect 1086 428 1090 432
rect 1118 738 1122 742
rect 1150 278 1154 282
rect 1118 268 1122 272
rect 1206 548 1210 552
rect 1166 278 1170 282
rect 1158 258 1162 262
rect 1246 868 1250 872
rect 1294 868 1298 872
rect 1238 528 1242 532
rect 1094 188 1098 192
rect 934 168 938 172
rect 1002 103 1006 107
rect 1009 103 1010 107
rect 1010 103 1013 107
rect 902 78 906 82
rect 1222 168 1226 172
rect 1286 468 1290 472
rect 1270 168 1274 172
rect 1334 548 1338 552
rect 1334 188 1338 192
rect 1270 78 1274 82
rect 942 48 946 52
rect 1310 48 1314 52
rect 482 3 486 7
rect 489 3 490 7
rect 490 3 493 7
<< metal5 >>
rect 1006 1303 1009 1307
rect 1005 1302 1010 1303
rect 1015 1302 1016 1307
rect 666 1268 742 1271
rect 486 1203 489 1207
rect 485 1202 490 1203
rect 495 1202 496 1207
rect 1006 1103 1009 1107
rect 1005 1102 1010 1103
rect 1015 1102 1016 1107
rect 338 1068 878 1071
rect 378 1058 462 1061
rect 322 1038 414 1041
rect 486 1003 489 1007
rect 485 1002 490 1003
rect 495 1002 496 1007
rect 1006 903 1009 907
rect 1005 902 1010 903
rect 1015 902 1016 907
rect 1250 868 1294 871
rect 330 848 406 851
rect 486 803 489 807
rect 485 802 490 803
rect 495 802 496 807
rect 194 738 230 741
rect 1010 738 1118 741
rect 1006 703 1009 707
rect 1005 702 1010 703
rect 1015 702 1016 707
rect 18 668 342 671
rect 818 668 1038 671
rect 1026 638 1070 641
rect 486 603 489 607
rect 485 602 490 603
rect 495 602 496 607
rect 978 558 1337 561
rect 1334 552 1337 558
rect 1010 548 1206 551
rect 802 528 1014 531
rect 1018 528 1238 531
rect 1006 503 1009 507
rect 1005 502 1010 503
rect 1015 502 1016 507
rect 514 478 702 481
rect 922 478 1054 481
rect 698 468 790 471
rect 986 468 1286 471
rect 402 458 446 461
rect 802 458 1006 461
rect 650 428 1086 431
rect 486 403 489 407
rect 485 402 490 403
rect 495 402 496 407
rect 34 348 94 351
rect 714 348 854 351
rect 1006 303 1009 307
rect 1005 302 1010 303
rect 1015 302 1016 307
rect 858 278 974 281
rect 978 278 1150 281
rect 922 268 942 271
rect 1166 271 1169 278
rect 1122 268 1169 271
rect 586 258 1158 261
rect 486 203 489 207
rect 485 202 490 203
rect 495 202 496 207
rect 1098 188 1334 191
rect 938 168 1222 171
rect 1226 168 1270 171
rect 1006 103 1009 107
rect 1005 102 1010 103
rect 1015 102 1016 107
rect 906 78 1270 81
rect 946 48 1310 51
rect 486 3 489 7
rect 485 2 490 3
rect 495 2 496 7
<< m6contact >>
rect 1000 1303 1002 1307
rect 1002 1303 1005 1307
rect 1010 1303 1013 1307
rect 1013 1303 1015 1307
rect 1000 1302 1005 1303
rect 1010 1302 1015 1303
rect 480 1203 482 1207
rect 482 1203 485 1207
rect 490 1203 493 1207
rect 493 1203 495 1207
rect 480 1202 485 1203
rect 490 1202 495 1203
rect 1000 1103 1002 1107
rect 1002 1103 1005 1107
rect 1010 1103 1013 1107
rect 1013 1103 1015 1107
rect 1000 1102 1005 1103
rect 1010 1102 1015 1103
rect 480 1003 482 1007
rect 482 1003 485 1007
rect 490 1003 493 1007
rect 493 1003 495 1007
rect 480 1002 485 1003
rect 490 1002 495 1003
rect 1000 903 1002 907
rect 1002 903 1005 907
rect 1010 903 1013 907
rect 1013 903 1015 907
rect 1000 902 1005 903
rect 1010 902 1015 903
rect 480 803 482 807
rect 482 803 485 807
rect 490 803 493 807
rect 493 803 495 807
rect 480 802 485 803
rect 490 802 495 803
rect 1000 703 1002 707
rect 1002 703 1005 707
rect 1010 703 1013 707
rect 1013 703 1015 707
rect 1000 702 1005 703
rect 1010 702 1015 703
rect 480 603 482 607
rect 482 603 485 607
rect 490 603 493 607
rect 493 603 495 607
rect 480 602 485 603
rect 490 602 495 603
rect 1000 503 1002 507
rect 1002 503 1005 507
rect 1010 503 1013 507
rect 1013 503 1015 507
rect 1000 502 1005 503
rect 1010 502 1015 503
rect 480 403 482 407
rect 482 403 485 407
rect 490 403 493 407
rect 493 403 495 407
rect 480 402 485 403
rect 490 402 495 403
rect 1000 303 1002 307
rect 1002 303 1005 307
rect 1010 303 1013 307
rect 1013 303 1015 307
rect 1000 302 1005 303
rect 1010 302 1015 303
rect 480 203 482 207
rect 482 203 485 207
rect 490 203 493 207
rect 493 203 495 207
rect 480 202 485 203
rect 490 202 495 203
rect 1000 103 1002 107
rect 1002 103 1005 107
rect 1010 103 1013 107
rect 1013 103 1015 107
rect 1000 102 1005 103
rect 1010 102 1015 103
rect 480 3 482 7
rect 482 3 485 7
rect 490 3 493 7
rect 493 3 495 7
rect 480 2 485 3
rect 490 2 495 3
<< metal6 >>
rect 480 1207 496 1330
rect 485 1202 490 1207
rect 495 1202 496 1207
rect 480 1007 496 1202
rect 485 1002 490 1007
rect 495 1002 496 1007
rect 480 807 496 1002
rect 485 802 490 807
rect 495 802 496 807
rect 480 607 496 802
rect 485 602 490 607
rect 495 602 496 607
rect 480 407 496 602
rect 485 402 490 407
rect 495 402 496 407
rect 480 207 496 402
rect 485 202 490 207
rect 495 202 496 207
rect 480 7 496 202
rect 485 2 490 7
rect 495 2 496 7
rect 480 -30 496 2
rect 1000 1307 1016 1330
rect 1005 1302 1010 1307
rect 1015 1302 1016 1307
rect 1000 1107 1016 1302
rect 1005 1102 1010 1107
rect 1015 1102 1016 1107
rect 1000 907 1016 1102
rect 1005 902 1010 907
rect 1015 902 1016 907
rect 1000 707 1016 902
rect 1005 702 1010 707
rect 1015 702 1016 707
rect 1000 507 1016 702
rect 1005 502 1010 507
rect 1015 502 1016 507
rect 1000 307 1016 502
rect 1005 302 1010 307
rect 1015 302 1016 307
rect 1000 107 1016 302
rect 1005 102 1010 107
rect 1015 102 1016 107
rect 1000 -30 1016 102
use OAI21X1  OAI21X1_17
timestamp 1751429576
transform -1 0 100 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_11
timestamp 1751429576
transform -1 0 68 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_12
timestamp 1751429576
transform -1 0 36 0 1 105
box -2 -3 34 103
use XOR2X1  XOR2X1_2
timestamp 1751429576
transform 1 0 60 0 -1 105
box -2 -3 58 103
use XNOR2X1  XNOR2X1_3
timestamp 1751429576
transform 1 0 4 0 -1 105
box -2 -3 58 103
use OAI21X1  OAI21X1_16
timestamp 1751429576
transform -1 0 164 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_10
timestamp 1751429576
transform -1 0 132 0 1 105
box -2 -3 34 103
use NOR3X1  NOR3X1_3
timestamp 1751429576
transform -1 0 180 0 -1 105
box -2 -3 66 103
use OAI21X1  OAI21X1_14
timestamp 1751429576
transform 1 0 164 0 1 105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_2
timestamp 1751429576
transform -1 0 236 0 -1 105
box -2 -3 58 103
use NAND3X1  NAND3X1_8
timestamp 1751429576
transform 1 0 228 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_9
timestamp 1751429576
transform -1 0 228 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_15
timestamp 1751429576
transform -1 0 284 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_6
timestamp 1751429576
transform 1 0 236 0 -1 105
box -2 -3 18 103
use AND2X2  AND2X2_3
timestamp 1751429576
transform 1 0 316 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_6
timestamp 1751429576
transform 1 0 292 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_8
timestamp 1751429576
transform -1 0 292 0 1 105
box -2 -3 34 103
use XOR2X1  XOR2X1_1
timestamp 1751429576
transform 1 0 284 0 -1 105
box -2 -3 58 103
use NAND3X1  NAND3X1_7
timestamp 1751429576
transform -1 0 380 0 1 105
box -2 -3 34 103
use NOR3X1  NOR3X1_2
timestamp 1751429576
transform 1 0 340 0 -1 105
box -2 -3 66 103
use BUFX4  BUFX4_13
timestamp 1751429576
transform 1 0 428 0 1 105
box -2 -3 34 103
use INVX1  INVX1_7
timestamp 1751429576
transform 1 0 412 0 1 105
box -2 -3 18 103
use AOI21X1  AOI21X1_7
timestamp 1751429576
transform -1 0 412 0 1 105
box -2 -3 34 103
use NOR3X1  NOR3X1_1
timestamp 1751429576
transform -1 0 468 0 -1 105
box -2 -3 66 103
use FILL  FILL_1_0_1
timestamp 1751429576
transform 1 0 500 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_0
timestamp 1751429576
transform 1 0 492 0 1 105
box -2 -3 10 103
use AOI21X1  AOI21X1_5
timestamp 1751429576
transform -1 0 492 0 1 105
box -2 -3 34 103
use FILL  FILL_0_0_0
timestamp 1751429576
transform -1 0 508 0 -1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_13
timestamp 1751429576
transform 1 0 468 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_3
timestamp 1751429576
transform 1 0 540 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_6
timestamp 1751429576
transform 1 0 508 0 1 105
box -2 -3 34 103
use BUFX4  BUFX4_6
timestamp 1751429576
transform 1 0 540 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_8
timestamp 1751429576
transform -1 0 540 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_0_1
timestamp 1751429576
transform -1 0 516 0 -1 105
box -2 -3 10 103
use MUX2X1  MUX2X1_4
timestamp 1751429576
transform -1 0 620 0 1 105
box -2 -3 50 103
use BUFX4  BUFX4_1
timestamp 1751429576
transform 1 0 596 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_1
timestamp 1751429576
transform 1 0 572 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_9
timestamp 1751429576
transform -1 0 660 0 1 105
box -2 -3 26 103
use INVX1  INVX1_39
timestamp 1751429576
transform 1 0 620 0 1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_63
timestamp 1751429576
transform 1 0 652 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_16
timestamp 1751429576
transform 1 0 628 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_1
timestamp 1751429576
transform 1 0 700 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_62
timestamp 1751429576
transform -1 0 700 0 1 105
box -2 -3 26 103
use INVX2  INVX2_22
timestamp 1751429576
transform 1 0 660 0 1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_73
timestamp 1751429576
transform 1 0 692 0 -1 105
box -2 -3 26 103
use INVX2  INVX2_4
timestamp 1751429576
transform 1 0 676 0 -1 105
box -2 -3 18 103
use INVX2  INVX2_24
timestamp 1751429576
transform -1 0 732 0 -1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_55
timestamp 1751429576
transform 1 0 780 0 1 105
box -2 -3 26 103
use INVX1  INVX1_1
timestamp 1751429576
transform 1 0 764 0 1 105
box -2 -3 18 103
use NAND3X1  NAND3X1_1
timestamp 1751429576
transform 1 0 732 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_24
timestamp 1751429576
transform 1 0 788 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_25
timestamp 1751429576
transform 1 0 756 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_1
timestamp 1751429576
transform 1 0 732 0 -1 105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_1
timestamp 1751429576
transform 1 0 804 0 1 105
box -2 -3 58 103
use INVX1  INVX1_3
timestamp 1751429576
transform 1 0 844 0 -1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_2
timestamp 1751429576
transform 1 0 820 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_2
timestamp 1751429576
transform 1 0 908 0 1 105
box -2 -3 34 103
use INVX2  INVX2_1
timestamp 1751429576
transform 1 0 892 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_3
timestamp 1751429576
transform -1 0 892 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_8
timestamp 1751429576
transform -1 0 916 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_6
timestamp 1751429576
transform -1 0 884 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_10
timestamp 1751429576
transform -1 0 972 0 1 105
box -2 -3 34 103
use OAI22X1  OAI22X1_2
timestamp 1751429576
transform -1 0 988 0 -1 105
box -2 -3 42 103
use OAI21X1  OAI21X1_27
timestamp 1751429576
transform -1 0 948 0 -1 105
box -2 -3 34 103
use AND2X2  AND2X2_2
timestamp 1751429576
transform -1 0 1004 0 1 105
box -2 -3 34 103
use FILL  FILL_0_1_1
timestamp 1751429576
transform 1 0 996 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_0
timestamp 1751429576
transform 1 0 988 0 -1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_59
timestamp 1751429576
transform 1 0 1020 0 1 105
box -2 -3 26 103
use FILL  FILL_1_1_1
timestamp 1751429576
transform 1 0 1012 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_0
timestamp 1751429576
transform 1 0 1004 0 1 105
box -2 -3 10 103
use INVX1  INVX1_37
timestamp 1751429576
transform -1 0 1052 0 -1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_93
timestamp 1751429576
transform 1 0 1004 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_2
timestamp 1751429576
transform 1 0 1076 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_5
timestamp 1751429576
transform 1 0 1044 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_4
timestamp 1751429576
transform 1 0 1084 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_4
timestamp 1751429576
transform 1 0 1052 0 -1 105
box -2 -3 34 103
use OAI22X1  OAI22X1_7
timestamp 1751429576
transform -1 0 1148 0 1 105
box -2 -3 42 103
use OAI22X1  OAI22X1_9
timestamp 1751429576
transform 1 0 1124 0 -1 105
box -2 -3 42 103
use INVX1  INVX1_41
timestamp 1751429576
transform 1 0 1108 0 -1 105
box -2 -3 18 103
use AND2X2  AND2X2_1
timestamp 1751429576
transform -1 0 1204 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_64
timestamp 1751429576
transform -1 0 1172 0 1 105
box -2 -3 26 103
use OR2X2  OR2X2_10
timestamp 1751429576
transform 1 0 1164 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_3
timestamp 1751429576
transform -1 0 1228 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_110
timestamp 1751429576
transform -1 0 1228 0 -1 105
box -2 -3 34 103
use INVX2  INVX2_23
timestamp 1751429576
transform 1 0 1268 0 1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_57
timestamp 1751429576
transform 1 0 1244 0 1 105
box -2 -3 26 103
use INVX2  INVX2_18
timestamp 1751429576
transform -1 0 1244 0 1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_14
timestamp 1751429576
transform 1 0 1252 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_12
timestamp 1751429576
transform 1 0 1228 0 -1 105
box -2 -3 26 103
use NAND3X1  NAND3X1_26
timestamp 1751429576
transform 1 0 1316 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_31
timestamp 1751429576
transform 1 0 1284 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_13
timestamp 1751429576
transform -1 0 1348 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_28
timestamp 1751429576
transform 1 0 1292 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_9
timestamp 1751429576
transform 1 0 1276 0 -1 105
box -2 -3 18 103
use OAI22X1  OAI22X1_5
timestamp 1751429576
transform -1 0 1412 0 1 105
box -2 -3 42 103
use NOR2X1  NOR2X1_16
timestamp 1751429576
transform 1 0 1348 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_21
timestamp 1751429576
transform 1 0 1396 0 -1 105
box -2 -3 34 103
use OR2X2  OR2X2_2
timestamp 1751429576
transform 1 0 1364 0 -1 105
box -2 -3 34 103
use INVX2  INVX2_3
timestamp 1751429576
transform 1 0 1348 0 -1 105
box -2 -3 18 103
use NOR3X1  NOR3X1_4
timestamp 1751429576
transform 1 0 1412 0 1 105
box -2 -3 66 103
use AOI21X1  AOI21X1_20
timestamp 1751429576
transform 1 0 1428 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_26
timestamp 1751429576
transform 1 0 1460 0 -1 105
box -2 -3 34 103
use FILL  FILL_1_1
timestamp 1751429576
transform -1 0 1500 0 -1 105
box -2 -3 10 103
use FILL  FILL_1_2
timestamp 1751429576
transform -1 0 1508 0 -1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_29
timestamp 1751429576
transform -1 0 1500 0 1 105
box -2 -3 26 103
use FILL  FILL_2_1
timestamp 1751429576
transform 1 0 1500 0 1 105
box -2 -3 10 103
use XNOR2X1  XNOR2X1_4
timestamp 1751429576
transform -1 0 60 0 -1 305
box -2 -3 58 103
use NAND3X1  NAND3X1_15
timestamp 1751429576
transform -1 0 92 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_15
timestamp 1751429576
transform 1 0 92 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_8
timestamp 1751429576
transform 1 0 124 0 -1 305
box -2 -3 18 103
use AOI21X1  AOI21X1_14
timestamp 1751429576
transform -1 0 172 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_16
timestamp 1751429576
transform 1 0 172 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_2
timestamp 1751429576
transform 1 0 204 0 -1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_4
timestamp 1751429576
transform -1 0 260 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_3
timestamp 1751429576
transform -1 0 292 0 -1 305
box -2 -3 34 103
use BUFX4  BUFX4_11
timestamp 1751429576
transform -1 0 324 0 -1 305
box -2 -3 34 103
use BUFX4  BUFX4_12
timestamp 1751429576
transform 1 0 324 0 -1 305
box -2 -3 34 103
use OAI22X1  OAI22X1_4
timestamp 1751429576
transform -1 0 396 0 -1 305
box -2 -3 42 103
use NAND3X1  NAND3X1_6
timestamp 1751429576
transform -1 0 428 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_5
timestamp 1751429576
transform 1 0 428 0 -1 305
box -2 -3 34 103
use BUFX4  BUFX4_2
timestamp 1751429576
transform -1 0 492 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_0_0
timestamp 1751429576
transform -1 0 500 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1751429576
transform -1 0 508 0 -1 305
box -2 -3 10 103
use INVX4  INVX4_2
timestamp 1751429576
transform -1 0 532 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_23
timestamp 1751429576
transform 1 0 532 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_41
timestamp 1751429576
transform -1 0 588 0 -1 305
box -2 -3 34 103
use AND2X2  AND2X2_5
timestamp 1751429576
transform -1 0 620 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_20
timestamp 1751429576
transform 1 0 620 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_44
timestamp 1751429576
transform -1 0 660 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_33
timestamp 1751429576
transform -1 0 692 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_32
timestamp 1751429576
transform 1 0 692 0 -1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_1
timestamp 1751429576
transform -1 0 764 0 -1 305
box -2 -3 50 103
use NOR2X1  NOR2X1_54
timestamp 1751429576
transform -1 0 788 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_14
timestamp 1751429576
transform 1 0 788 0 -1 305
box -2 -3 18 103
use AOI21X1  AOI21X1_39
timestamp 1751429576
transform 1 0 804 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_105
timestamp 1751429576
transform 1 0 836 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_9
timestamp 1751429576
transform -1 0 900 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_2
timestamp 1751429576
transform -1 0 916 0 -1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_58
timestamp 1751429576
transform -1 0 940 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_32
timestamp 1751429576
transform 1 0 940 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_51
timestamp 1751429576
transform 1 0 972 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_1_0
timestamp 1751429576
transform 1 0 996 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1751429576
transform 1 0 1004 0 -1 305
box -2 -3 10 103
use AND2X2  AND2X2_11
timestamp 1751429576
transform 1 0 1012 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_35
timestamp 1751429576
transform -1 0 1060 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_87
timestamp 1751429576
transform -1 0 1092 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_52
timestamp 1751429576
transform 1 0 1092 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_50
timestamp 1751429576
transform 1 0 1124 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_64
timestamp 1751429576
transform 1 0 1156 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_94
timestamp 1751429576
transform -1 0 1220 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_89
timestamp 1751429576
transform -1 0 1252 0 -1 305
box -2 -3 34 103
use AND2X2  AND2X2_10
timestamp 1751429576
transform 1 0 1252 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_60
timestamp 1751429576
transform 1 0 1284 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_65
timestamp 1751429576
transform -1 0 1332 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_106
timestamp 1751429576
transform 1 0 1332 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_63
timestamp 1751429576
transform 1 0 1364 0 -1 305
box -2 -3 34 103
use INVX4  INVX4_3
timestamp 1751429576
transform -1 0 1420 0 -1 305
box -2 -3 26 103
use INVX2  INVX2_8
timestamp 1751429576
transform -1 0 1436 0 -1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_30
timestamp 1751429576
transform 1 0 1436 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_22
timestamp 1751429576
transform -1 0 1484 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_17
timestamp 1751429576
transform 1 0 1484 0 -1 305
box -2 -3 18 103
use FILL  FILL_3_1
timestamp 1751429576
transform -1 0 1508 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_19
timestamp 1751429576
transform -1 0 36 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_11
timestamp 1751429576
transform 1 0 36 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_13
timestamp 1751429576
transform 1 0 68 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_21
timestamp 1751429576
transform 1 0 100 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_17
timestamp 1751429576
transform 1 0 132 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_12
timestamp 1751429576
transform -1 0 196 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_10
timestamp 1751429576
transform 1 0 196 0 1 305
box -2 -3 34 103
use XOR2X1  XOR2X1_3
timestamp 1751429576
transform 1 0 228 0 1 305
box -2 -3 58 103
use NAND2X1  NAND2X1_5
timestamp 1751429576
transform -1 0 308 0 1 305
box -2 -3 26 103
use INVX1  INVX1_43
timestamp 1751429576
transform -1 0 324 0 1 305
box -2 -3 18 103
use BUFX4  BUFX4_10
timestamp 1751429576
transform 1 0 324 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_66
timestamp 1751429576
transform -1 0 380 0 1 305
box -2 -3 26 103
use BUFX4  BUFX4_14
timestamp 1751429576
transform 1 0 380 0 1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_10
timestamp 1751429576
transform -1 0 452 0 1 305
box -2 -3 42 103
use NAND2X1  NAND2X1_7
timestamp 1751429576
transform -1 0 476 0 1 305
box -2 -3 26 103
use FILL  FILL_3_0_0
timestamp 1751429576
transform -1 0 484 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1751429576
transform -1 0 492 0 1 305
box -2 -3 10 103
use BUFX4  BUFX4_9
timestamp 1751429576
transform -1 0 524 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_7
timestamp 1751429576
transform 1 0 524 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_8
timestamp 1751429576
transform 1 0 556 0 1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_5
timestamp 1751429576
transform 1 0 588 0 1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_3
timestamp 1751429576
transform -1 0 684 0 1 305
box -2 -3 50 103
use OAI21X1  OAI21X1_107
timestamp 1751429576
transform 1 0 684 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_27
timestamp 1751429576
transform 1 0 716 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_6
timestamp 1751429576
transform 1 0 748 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_32
timestamp 1751429576
transform -1 0 812 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_29
timestamp 1751429576
transform 1 0 812 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_31
timestamp 1751429576
transform -1 0 868 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_15
timestamp 1751429576
transform 1 0 868 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_22
timestamp 1751429576
transform -1 0 924 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_14
timestamp 1751429576
transform -1 0 948 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_30
timestamp 1751429576
transform 1 0 948 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_1
timestamp 1751429576
transform -1 0 1012 0 1 305
box -2 -3 34 103
use FILL  FILL_3_1_0
timestamp 1751429576
transform -1 0 1020 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1751429576
transform -1 0 1028 0 1 305
box -2 -3 10 103
use NAND2X1  NAND2X1_61
timestamp 1751429576
transform -1 0 1052 0 1 305
box -2 -3 26 103
use INVX2  INVX2_9
timestamp 1751429576
transform -1 0 1068 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_108
timestamp 1751429576
transform -1 0 1100 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_66
timestamp 1751429576
transform -1 0 1124 0 1 305
box -2 -3 26 103
use AND2X2  AND2X2_12
timestamp 1751429576
transform 1 0 1124 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_111
timestamp 1751429576
transform 1 0 1156 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_59
timestamp 1751429576
transform 1 0 1188 0 1 305
box -2 -3 26 103
use OR2X2  OR2X2_9
timestamp 1751429576
transform 1 0 1212 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_62
timestamp 1751429576
transform 1 0 1244 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_67
timestamp 1751429576
transform 1 0 1276 0 1 305
box -2 -3 26 103
use OR2X2  OR2X2_11
timestamp 1751429576
transform -1 0 1332 0 1 305
box -2 -3 34 103
use INVX2  INVX2_11
timestamp 1751429576
transform -1 0 1348 0 1 305
box -2 -3 18 103
use NAND3X1  NAND3X1_29
timestamp 1751429576
transform -1 0 1380 0 1 305
box -2 -3 34 103
use OR2X2  OR2X2_4
timestamp 1751429576
transform -1 0 1412 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_33
timestamp 1751429576
transform -1 0 1436 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_20
timestamp 1751429576
transform -1 0 1460 0 1 305
box -2 -3 26 103
use OR2X2  OR2X2_3
timestamp 1751429576
transform -1 0 1492 0 1 305
box -2 -3 34 103
use FILL  FILL_4_1
timestamp 1751429576
transform 1 0 1492 0 1 305
box -2 -3 10 103
use FILL  FILL_4_2
timestamp 1751429576
transform 1 0 1500 0 1 305
box -2 -3 10 103
use AND2X2  AND2X2_4
timestamp 1751429576
transform -1 0 36 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_4
timestamp 1751429576
transform 1 0 36 0 -1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_14
timestamp 1751429576
transform -1 0 92 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_3
timestamp 1751429576
transform 1 0 92 0 -1 505
box -2 -3 26 103
use INVX1  INVX1_5
timestamp 1751429576
transform 1 0 116 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_12
timestamp 1751429576
transform 1 0 132 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_8
timestamp 1751429576
transform -1 0 188 0 -1 505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_5
timestamp 1751429576
transform -1 0 244 0 -1 505
box -2 -3 58 103
use AOI21X1  AOI21X1_74
timestamp 1751429576
transform -1 0 276 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_120
timestamp 1751429576
transform -1 0 308 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_117
timestamp 1751429576
transform -1 0 340 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_121
timestamp 1751429576
transform 1 0 340 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_118
timestamp 1751429576
transform -1 0 404 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_71
timestamp 1751429576
transform -1 0 428 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_68
timestamp 1751429576
transform -1 0 460 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_65
timestamp 1751429576
transform -1 0 484 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_0_0
timestamp 1751429576
transform -1 0 492 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1751429576
transform -1 0 500 0 -1 505
box -2 -3 10 103
use AOI21X1  AOI21X1_69
timestamp 1751429576
transform -1 0 532 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_57
timestamp 1751429576
transform -1 0 556 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_56
timestamp 1751429576
transform 1 0 556 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_119
timestamp 1751429576
transform -1 0 612 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_15
timestamp 1751429576
transform -1 0 636 0 -1 505
box -2 -3 26 103
use BUFX4  BUFX4_4
timestamp 1751429576
transform -1 0 668 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_5
timestamp 1751429576
transform 1 0 668 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_48
timestamp 1751429576
transform -1 0 724 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_67
timestamp 1751429576
transform -1 0 748 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_40
timestamp 1751429576
transform -1 0 780 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_5
timestamp 1751429576
transform -1 0 804 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_71
timestamp 1751429576
transform 1 0 804 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_90
timestamp 1751429576
transform 1 0 836 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_60
timestamp 1751429576
transform -1 0 900 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_91
timestamp 1751429576
transform 1 0 900 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_50
timestamp 1751429576
transform -1 0 956 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_7
timestamp 1751429576
transform 1 0 956 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_1_0
timestamp 1751429576
transform -1 0 996 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1751429576
transform -1 0 1004 0 -1 505
box -2 -3 10 103
use OAI22X1  OAI22X1_1
timestamp 1751429576
transform -1 0 1044 0 -1 505
box -2 -3 42 103
use OAI21X1  OAI21X1_61
timestamp 1751429576
transform -1 0 1076 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_92
timestamp 1751429576
transform 1 0 1076 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_40
timestamp 1751429576
transform -1 0 1124 0 -1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_40
timestamp 1751429576
transform 1 0 1124 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_109
timestamp 1751429576
transform 1 0 1148 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_73
timestamp 1751429576
transform 1 0 1180 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_24
timestamp 1751429576
transform -1 0 1236 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_28
timestamp 1751429576
transform 1 0 1236 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_38
timestamp 1751429576
transform -1 0 1300 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_25
timestamp 1751429576
transform 1 0 1300 0 -1 505
box -2 -3 34 103
use INVX2  INVX2_7
timestamp 1751429576
transform -1 0 1348 0 -1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_28
timestamp 1751429576
transform 1 0 1348 0 -1 505
box -2 -3 26 103
use INVX4  INVX4_7
timestamp 1751429576
transform -1 0 1396 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_25
timestamp 1751429576
transform 1 0 1396 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_21
timestamp 1751429576
transform -1 0 1452 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_37
timestamp 1751429576
transform -1 0 1484 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_31
timestamp 1751429576
transform 1 0 1484 0 -1 505
box -2 -3 26 103
use INVX1  INVX1_4
timestamp 1751429576
transform 1 0 4 0 1 505
box -2 -3 18 103
use NAND3X1  NAND3X1_2
timestamp 1751429576
transform 1 0 20 0 1 505
box -2 -3 34 103
use OR2X2  OR2X2_1
timestamp 1751429576
transform -1 0 84 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_18
timestamp 1751429576
transform -1 0 116 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_124
timestamp 1751429576
transform -1 0 148 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_9
timestamp 1751429576
transform 1 0 148 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_67
timestamp 1751429576
transform 1 0 180 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_68
timestamp 1751429576
transform -1 0 244 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_66
timestamp 1751429576
transform -1 0 276 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_73
timestamp 1751429576
transform -1 0 308 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_65
timestamp 1751429576
transform 1 0 308 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_69
timestamp 1751429576
transform 1 0 340 0 1 505
box -2 -3 34 103
use OAI22X1  OAI22X1_10
timestamp 1751429576
transform 1 0 372 0 1 505
box -2 -3 42 103
use AOI22X1  AOI22X1_8
timestamp 1751429576
transform -1 0 452 0 1 505
box -2 -3 42 103
use AOI21X1  AOI21X1_70
timestamp 1751429576
transform -1 0 484 0 1 505
box -2 -3 34 103
use FILL  FILL_5_0_0
timestamp 1751429576
transform -1 0 492 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1751429576
transform -1 0 500 0 1 505
box -2 -3 10 103
use INVX2  INVX2_20
timestamp 1751429576
transform -1 0 516 0 1 505
box -2 -3 18 103
use AOI21X1  AOI21X1_57
timestamp 1751429576
transform -1 0 548 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_61
timestamp 1751429576
transform 1 0 548 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_56
timestamp 1751429576
transform -1 0 604 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_37
timestamp 1751429576
transform 1 0 604 0 1 505
box -2 -3 26 103
use INVX8  INVX8_2
timestamp 1751429576
transform 1 0 628 0 1 505
box -2 -3 42 103
use NOR2X1  NOR2X1_7
timestamp 1751429576
transform 1 0 668 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_24
timestamp 1751429576
transform 1 0 692 0 1 505
box -2 -3 26 103
use INVX1  INVX1_15
timestamp 1751429576
transform -1 0 732 0 1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_23
timestamp 1751429576
transform -1 0 756 0 1 505
box -2 -3 26 103
use INVX2  INVX2_17
timestamp 1751429576
transform -1 0 772 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_56
timestamp 1751429576
transform -1 0 804 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_17
timestamp 1751429576
transform 1 0 804 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_27
timestamp 1751429576
transform -1 0 852 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_57
timestamp 1751429576
transform 1 0 852 0 1 505
box -2 -3 34 103
use INVX1  INVX1_36
timestamp 1751429576
transform 1 0 884 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_58
timestamp 1751429576
transform 1 0 900 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_35
timestamp 1751429576
transform 1 0 932 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_25
timestamp 1751429576
transform 1 0 964 0 1 505
box -2 -3 26 103
use FILL  FILL_5_1_0
timestamp 1751429576
transform 1 0 988 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1751429576
transform 1 0 996 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_34
timestamp 1751429576
transform 1 0 1004 0 1 505
box -2 -3 34 103
use INVX1  INVX1_16
timestamp 1751429576
transform 1 0 1036 0 1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_34
timestamp 1751429576
transform 1 0 1052 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_51
timestamp 1751429576
transform -1 0 1108 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_46
timestamp 1751429576
transform 1 0 1108 0 1 505
box -2 -3 34 103
use INVX1  INVX1_22
timestamp 1751429576
transform 1 0 1140 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_36
timestamp 1751429576
transform 1 0 1156 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_45
timestamp 1751429576
transform 1 0 1188 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_26
timestamp 1751429576
transform -1 0 1236 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_24
timestamp 1751429576
transform 1 0 1236 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_74
timestamp 1751429576
transform 1 0 1268 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_40
timestamp 1751429576
transform -1 0 1332 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_37
timestamp 1751429576
transform 1 0 1332 0 1 505
box -2 -3 34 103
use INVX4  INVX4_5
timestamp 1751429576
transform 1 0 1364 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_47
timestamp 1751429576
transform 1 0 1388 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_35
timestamp 1751429576
transform 1 0 1420 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_39
timestamp 1751429576
transform -1 0 1468 0 1 505
box -2 -3 26 103
use INVX1  INVX1_18
timestamp 1751429576
transform -1 0 1484 0 1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_32
timestamp 1751429576
transform 1 0 1484 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_13
timestamp 1751429576
transform 1 0 4 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_10
timestamp 1751429576
transform 1 0 36 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_16
timestamp 1751429576
transform -1 0 92 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_18
timestamp 1751429576
transform 1 0 92 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_72
timestamp 1751429576
transform -1 0 156 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_70
timestamp 1751429576
transform 1 0 156 0 -1 705
box -2 -3 34 103
use AND2X2  AND2X2_13
timestamp 1751429576
transform -1 0 220 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_70
timestamp 1751429576
transform -1 0 244 0 -1 705
box -2 -3 26 103
use OAI22X1  OAI22X1_3
timestamp 1751429576
transform -1 0 284 0 -1 705
box -2 -3 42 103
use NAND2X1  NAND2X1_40
timestamp 1751429576
transform -1 0 308 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_66
timestamp 1751429576
transform -1 0 340 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_54
timestamp 1751429576
transform -1 0 364 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_63
timestamp 1751429576
transform -1 0 388 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_99
timestamp 1751429576
transform -1 0 420 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_96
timestamp 1751429576
transform 1 0 420 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_98
timestamp 1751429576
transform -1 0 484 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_0_0
timestamp 1751429576
transform 1 0 484 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1751429576
transform 1 0 492 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_97
timestamp 1751429576
transform 1 0 500 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_53
timestamp 1751429576
transform -1 0 556 0 -1 705
box -2 -3 26 103
use OAI22X1  OAI22X1_8
timestamp 1751429576
transform 1 0 556 0 -1 705
box -2 -3 42 103
use AOI22X1  AOI22X1_6
timestamp 1751429576
transform -1 0 636 0 -1 705
box -2 -3 42 103
use AOI21X1  AOI21X1_45
timestamp 1751429576
transform -1 0 668 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_44
timestamp 1751429576
transform 1 0 668 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_39
timestamp 1751429576
transform 1 0 700 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_30
timestamp 1751429576
transform -1 0 748 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_39
timestamp 1751429576
transform 1 0 748 0 -1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_2
timestamp 1751429576
transform 1 0 780 0 -1 705
box -2 -3 50 103
use NAND2X1  NAND2X1_25
timestamp 1751429576
transform 1 0 828 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_18
timestamp 1751429576
transform 1 0 852 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_49
timestamp 1751429576
transform 1 0 876 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_31
timestamp 1751429576
transform 1 0 900 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_72
timestamp 1751429576
transform 1 0 916 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_56
timestamp 1751429576
transform 1 0 948 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_41
timestamp 1751429576
transform -1 0 996 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_1_0
timestamp 1751429576
transform 1 0 996 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1751429576
transform 1 0 1004 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_62
timestamp 1751429576
transform 1 0 1012 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_26
timestamp 1751429576
transform 1 0 1044 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_86
timestamp 1751429576
transform -1 0 1100 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_85
timestamp 1751429576
transform -1 0 1132 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_46
timestamp 1751429576
transform -1 0 1156 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_63
timestamp 1751429576
transform 1 0 1156 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_42
timestamp 1751429576
transform 1 0 1188 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_33
timestamp 1751429576
transform 1 0 1212 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_88
timestamp 1751429576
transform -1 0 1268 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_29
timestamp 1751429576
transform 1 0 1268 0 -1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_41
timestamp 1751429576
transform 1 0 1284 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_23
timestamp 1751429576
transform 1 0 1308 0 -1 705
box -2 -3 18 103
use AOI22X1  AOI22X1_4
timestamp 1751429576
transform 1 0 1324 0 -1 705
box -2 -3 42 103
use AOI22X1  AOI22X1_3
timestamp 1751429576
transform -1 0 1404 0 -1 705
box -2 -3 42 103
use NAND3X1  NAND3X1_30
timestamp 1751429576
transform 1 0 1404 0 -1 705
box -2 -3 34 103
use OR2X2  OR2X2_7
timestamp 1751429576
transform -1 0 1468 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_38
timestamp 1751429576
transform -1 0 1500 0 -1 705
box -2 -3 34 103
use FILL  FILL_7_1
timestamp 1751429576
transform -1 0 1508 0 -1 705
box -2 -3 10 103
use NAND3X1  NAND3X1_19
timestamp 1751429576
transform -1 0 36 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_20
timestamp 1751429576
transform -1 0 68 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_75
timestamp 1751429576
transform -1 0 100 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_77
timestamp 1751429576
transform -1 0 132 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_73
timestamp 1751429576
transform 1 0 132 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_68
timestamp 1751429576
transform -1 0 188 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_123
timestamp 1751429576
transform 1 0 188 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_115
timestamp 1751429576
transform 1 0 220 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_64
timestamp 1751429576
transform -1 0 276 0 1 705
box -2 -3 26 103
use INVX1  INVX1_42
timestamp 1751429576
transform 1 0 276 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_122
timestamp 1751429576
transform -1 0 324 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_116
timestamp 1751429576
transform 1 0 324 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_62
timestamp 1751429576
transform -1 0 380 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_67
timestamp 1751429576
transform -1 0 412 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_43
timestamp 1751429576
transform -1 0 444 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_55
timestamp 1751429576
transform -1 0 476 0 1 705
box -2 -3 34 103
use FILL  FILL_7_0_0
timestamp 1751429576
transform 1 0 476 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1751429576
transform 1 0 484 0 1 705
box -2 -3 10 103
use NAND3X1  NAND3X1_45
timestamp 1751429576
transform 1 0 492 0 1 705
box -2 -3 34 103
use INVX1  INVX1_38
timestamp 1751429576
transform -1 0 540 0 1 705
box -2 -3 18 103
use NAND3X1  NAND3X1_49
timestamp 1751429576
transform 1 0 540 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_44
timestamp 1751429576
transform 1 0 572 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_69
timestamp 1751429576
transform -1 0 628 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_78
timestamp 1751429576
transform -1 0 660 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_80
timestamp 1751429576
transform 1 0 660 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_52
timestamp 1751429576
transform 1 0 692 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_77
timestamp 1751429576
transform 1 0 716 0 1 705
box -2 -3 34 103
use INVX2  INVX2_12
timestamp 1751429576
transform 1 0 748 0 1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_22
timestamp 1751429576
transform 1 0 764 0 1 705
box -2 -3 26 103
use INVX4  INVX4_6
timestamp 1751429576
transform 1 0 788 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_29
timestamp 1751429576
transform 1 0 812 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_53
timestamp 1751429576
transform 1 0 836 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_51
timestamp 1751429576
transform -1 0 892 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_45
timestamp 1751429576
transform 1 0 892 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_28
timestamp 1751429576
transform 1 0 924 0 1 705
box -2 -3 26 103
use AND2X2  AND2X2_8
timestamp 1751429576
transform 1 0 948 0 1 705
box -2 -3 34 103
use AOI22X1  AOI22X1_2
timestamp 1751429576
transform -1 0 1020 0 1 705
box -2 -3 42 103
use FILL  FILL_7_1_0
timestamp 1751429576
transform -1 0 1028 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1751429576
transform -1 0 1036 0 1 705
box -2 -3 10 103
use INVX1  INVX1_24
timestamp 1751429576
transform -1 0 1052 0 1 705
box -2 -3 18 103
use AOI21X1  AOI21X1_49
timestamp 1751429576
transform -1 0 1084 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_30
timestamp 1751429576
transform 1 0 1084 0 1 705
box -2 -3 34 103
use AND2X2  AND2X2_7
timestamp 1751429576
transform -1 0 1148 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_37
timestamp 1751429576
transform -1 0 1172 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_43
timestamp 1751429576
transform -1 0 1204 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_27
timestamp 1751429576
transform -1 0 1228 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_37
timestamp 1751429576
transform -1 0 1260 0 1 705
box -2 -3 34 103
use AND2X2  AND2X2_6
timestamp 1751429576
transform 1 0 1260 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_36
timestamp 1751429576
transform -1 0 1316 0 1 705
box -2 -3 26 103
use INVX2  INVX2_6
timestamp 1751429576
transform 1 0 1316 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_44
timestamp 1751429576
transform 1 0 1332 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_42
timestamp 1751429576
transform 1 0 1364 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_48
timestamp 1751429576
transform -1 0 1428 0 1 705
box -2 -3 34 103
use OR2X2  OR2X2_5
timestamp 1751429576
transform 1 0 1428 0 1 705
box -2 -3 34 103
use INVX2  INVX2_16
timestamp 1751429576
transform -1 0 1476 0 1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_42
timestamp 1751429576
transform 1 0 1476 0 1 705
box -2 -3 26 103
use FILL  FILL_8_1
timestamp 1751429576
transform 1 0 1500 0 1 705
box -2 -3 10 103
use AOI21X1  AOI21X1_4
timestamp 1751429576
transform 1 0 4 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_125
timestamp 1751429576
transform -1 0 68 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_76
timestamp 1751429576
transform -1 0 100 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_76
timestamp 1751429576
transform -1 0 132 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_74
timestamp 1751429576
transform -1 0 164 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_71
timestamp 1751429576
transform 1 0 164 0 -1 905
box -2 -3 34 103
use XOR2X1  XOR2X1_5
timestamp 1751429576
transform 1 0 196 0 -1 905
box -2 -3 58 103
use NAND2X1  NAND2X1_9
timestamp 1751429576
transform -1 0 276 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_113
timestamp 1751429576
transform -1 0 308 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_114
timestamp 1751429576
transform -1 0 340 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_50
timestamp 1751429576
transform -1 0 372 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_65
timestamp 1751429576
transform -1 0 404 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_47
timestamp 1751429576
transform -1 0 428 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_58
timestamp 1751429576
transform -1 0 452 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_100
timestamp 1751429576
transform -1 0 484 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_0_0
timestamp 1751429576
transform 1 0 484 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1751429576
transform 1 0 492 0 -1 905
box -2 -3 10 103
use NAND2X1  NAND2X1_55
timestamp 1751429576
transform 1 0 500 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_95
timestamp 1751429576
transform 1 0 524 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_54
timestamp 1751429576
transform 1 0 556 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_52
timestamp 1751429576
transform -1 0 612 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_46
timestamp 1751429576
transform -1 0 636 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_75
timestamp 1751429576
transform -1 0 668 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_79
timestamp 1751429576
transform -1 0 700 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_81
timestamp 1751429576
transform 1 0 700 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_35
timestamp 1751429576
transform -1 0 756 0 -1 905
box -2 -3 26 103
use XOR2X1  XOR2X1_4
timestamp 1751429576
transform -1 0 812 0 -1 905
box -2 -3 58 103
use AND2X2  AND2X2_9
timestamp 1751429576
transform 1 0 812 0 -1 905
box -2 -3 34 103
use INVX2  INVX2_10
timestamp 1751429576
transform -1 0 860 0 -1 905
box -2 -3 18 103
use INVX4  INVX4_4
timestamp 1751429576
transform 1 0 860 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_54
timestamp 1751429576
transform 1 0 884 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_33
timestamp 1751429576
transform -1 0 948 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_43
timestamp 1751429576
transform 1 0 948 0 -1 905
box -2 -3 26 103
use INVX1  INVX1_25
timestamp 1751429576
transform 1 0 972 0 -1 905
box -2 -3 18 103
use FILL  FILL_8_1_0
timestamp 1751429576
transform -1 0 996 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1751429576
transform -1 0 1004 0 -1 905
box -2 -3 10 103
use XNOR2X1  XNOR2X1_6
timestamp 1751429576
transform -1 0 1060 0 -1 905
box -2 -3 58 103
use NAND2X1  NAND2X1_36
timestamp 1751429576
transform -1 0 1084 0 -1 905
box -2 -3 26 103
use INVX4  INVX4_1
timestamp 1751429576
transform -1 0 1108 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_31
timestamp 1751429576
transform 1 0 1108 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_52
timestamp 1751429576
transform -1 0 1172 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_50
timestamp 1751429576
transform -1 0 1196 0 -1 905
box -2 -3 26 103
use OR2X2  OR2X2_6
timestamp 1751429576
transform 1 0 1196 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_29
timestamp 1751429576
transform 1 0 1228 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_51
timestamp 1751429576
transform 1 0 1260 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_50
timestamp 1751429576
transform 1 0 1292 0 -1 905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_7
timestamp 1751429576
transform 1 0 1324 0 -1 905
box -2 -3 58 103
use AOI21X1  AOI21X1_41
timestamp 1751429576
transform 1 0 1380 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_49
timestamp 1751429576
transform -1 0 1444 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_19
timestamp 1751429576
transform -1 0 1460 0 -1 905
box -2 -3 18 103
use BUFX2  BUFX2_1
timestamp 1751429576
transform 1 0 1460 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_43
timestamp 1751429576
transform -1 0 1508 0 -1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_79
timestamp 1751429576
transform -1 0 36 0 1 905
box -2 -3 34 103
use INVX2  INVX2_25
timestamp 1751429576
transform 1 0 36 0 1 905
box -2 -3 18 103
use NAND3X1  NAND3X1_77
timestamp 1751429576
transform -1 0 84 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_11
timestamp 1751429576
transform 1 0 84 0 1 905
box -2 -3 26 103
use AOI22X1  AOI22X1_1
timestamp 1751429576
transform 1 0 108 0 1 905
box -2 -3 42 103
use NAND3X1  NAND3X1_21
timestamp 1751429576
transform -1 0 180 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_19
timestamp 1751429576
transform 1 0 180 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_23
timestamp 1751429576
transform 1 0 212 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_72
timestamp 1751429576
transform -1 0 276 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_53
timestamp 1751429576
transform -1 0 308 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_52
timestamp 1751429576
transform -1 0 340 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_71
timestamp 1751429576
transform -1 0 372 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_51
timestamp 1751429576
transform 1 0 372 0 1 905
box -2 -3 34 103
use INVX2  INVX2_21
timestamp 1751429576
transform -1 0 420 0 1 905
box -2 -3 18 103
use NAND3X1  NAND3X1_47
timestamp 1751429576
transform 1 0 420 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_54
timestamp 1751429576
transform 1 0 452 0 1 905
box -2 -3 34 103
use FILL  FILL_9_0_0
timestamp 1751429576
transform 1 0 484 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1751429576
transform 1 0 492 0 1 905
box -2 -3 10 103
use NAND3X1  NAND3X1_48
timestamp 1751429576
transform 1 0 500 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_46
timestamp 1751429576
transform 1 0 532 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_60
timestamp 1751429576
transform -1 0 588 0 1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_39
timestamp 1751429576
transform -1 0 620 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_46
timestamp 1751429576
transform -1 0 652 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_47
timestamp 1751429576
transform -1 0 684 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_38
timestamp 1751429576
transform 1 0 684 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_43
timestamp 1751429576
transform -1 0 748 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_48
timestamp 1751429576
transform -1 0 772 0 1 905
box -2 -3 26 103
use OAI22X1  OAI22X1_6
timestamp 1751429576
transform 1 0 772 0 1 905
box -2 -3 42 103
use OAI21X1  OAI21X1_66
timestamp 1751429576
transform -1 0 844 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_67
timestamp 1751429576
transform 1 0 844 0 1 905
box -2 -3 34 103
use INVX2  INVX2_15
timestamp 1751429576
transform -1 0 892 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_68
timestamp 1751429576
transform -1 0 924 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_47
timestamp 1751429576
transform -1 0 948 0 1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_31
timestamp 1751429576
transform -1 0 980 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_55
timestamp 1751429576
transform 1 0 980 0 1 905
box -2 -3 34 103
use FILL  FILL_9_1_0
timestamp 1751429576
transform 1 0 1012 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1751429576
transform 1 0 1020 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_59
timestamp 1751429576
transform 1 0 1028 0 1 905
box -2 -3 34 103
use INVX1  INVX1_21
timestamp 1751429576
transform -1 0 1076 0 1 905
box -2 -3 18 103
use NOR2X1  NOR2X1_38
timestamp 1751429576
transform -1 0 1100 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_45
timestamp 1751429576
transform -1 0 1124 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_34
timestamp 1751429576
transform -1 0 1148 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_64
timestamp 1751429576
transform 1 0 1148 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_26
timestamp 1751429576
transform 1 0 1180 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_21
timestamp 1751429576
transform 1 0 1212 0 1 905
box -2 -3 26 103
use DFFSR  DFFSR_2
timestamp 1751429576
transform 1 0 1236 0 1 905
box -2 -3 178 103
use BUFX2  BUFX2_3
timestamp 1751429576
transform 1 0 1412 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_19
timestamp 1751429576
transform 1 0 1436 0 1 905
box -2 -3 26 103
use BUFX2  BUFX2_2
timestamp 1751429576
transform 1 0 1460 0 1 905
box -2 -3 26 103
use INVX1  INVX1_30
timestamp 1751429576
transform 1 0 1484 0 1 905
box -2 -3 18 103
use FILL  FILL_10_1
timestamp 1751429576
transform 1 0 1500 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_22
timestamp 1751429576
transform -1 0 36 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_17
timestamp 1751429576
transform -1 0 68 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_20
timestamp 1751429576
transform -1 0 100 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_23
timestamp 1751429576
transform 1 0 100 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_13
timestamp 1751429576
transform 1 0 132 0 -1 1105
box -2 -3 26 103
use INVX2  INVX2_2
timestamp 1751429576
transform 1 0 156 0 -1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_12
timestamp 1751429576
transform 1 0 172 0 -1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_22
timestamp 1751429576
transform -1 0 228 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_24
timestamp 1751429576
transform -1 0 260 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_59
timestamp 1751429576
transform -1 0 292 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_55
timestamp 1751429576
transform 1 0 292 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_60
timestamp 1751429576
transform 1 0 324 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_61
timestamp 1751429576
transform -1 0 388 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_58
timestamp 1751429576
transform -1 0 420 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_56
timestamp 1751429576
transform 1 0 420 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_59
timestamp 1751429576
transform 1 0 452 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_0_0
timestamp 1751429576
transform 1 0 484 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1751429576
transform 1 0 492 0 -1 1105
box -2 -3 10 103
use NAND3X1  NAND3X1_40
timestamp 1751429576
transform 1 0 500 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_101
timestamp 1751429576
transform -1 0 564 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_82
timestamp 1751429576
transform -1 0 596 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_48
timestamp 1751429576
transform 1 0 596 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_76
timestamp 1751429576
transform 1 0 628 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_83
timestamp 1751429576
transform -1 0 692 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_32
timestamp 1751429576
transform -1 0 724 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_36
timestamp 1751429576
transform -1 0 756 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_38
timestamp 1751429576
transform 1 0 756 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_27
timestamp 1751429576
transform -1 0 796 0 -1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_35
timestamp 1751429576
transform -1 0 828 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_33
timestamp 1751429576
transform 1 0 828 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_26
timestamp 1751429576
transform 1 0 860 0 -1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_23
timestamp 1751429576
transform 1 0 876 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_3
timestamp 1751429576
transform 1 0 908 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_68
timestamp 1751429576
transform -1 0 964 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_17
timestamp 1751429576
transform -1 0 988 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_44
timestamp 1751429576
transform 1 0 988 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_1_0
timestamp 1751429576
transform 1 0 1012 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1751429576
transform 1 0 1020 0 -1 1105
box -2 -3 10 103
use DFFSR  DFFSR_1
timestamp 1751429576
transform 1 0 1028 0 -1 1105
box -2 -3 178 103
use OAI21X1  OAI21X1_65
timestamp 1751429576
transform -1 0 1236 0 -1 1105
box -2 -3 34 103
use DFFSR  DFFSR_3
timestamp 1751429576
transform 1 0 1236 0 -1 1105
box -2 -3 178 103
use INVX1  INVX1_13
timestamp 1751429576
transform 1 0 1412 0 -1 1105
box -2 -3 18 103
use NAND3X1  NAND3X1_28
timestamp 1751429576
transform 1 0 1428 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_20
timestamp 1751429576
transform 1 0 1460 0 -1 1105
box -2 -3 26 103
use FILL  FILL_11_1
timestamp 1751429576
transform -1 0 1492 0 -1 1105
box -2 -3 10 103
use FILL  FILL_11_2
timestamp 1751429576
transform -1 0 1500 0 -1 1105
box -2 -3 10 103
use FILL  FILL_11_3
timestamp 1751429576
transform -1 0 1508 0 -1 1105
box -2 -3 10 103
use NAND3X1  NAND3X1_80
timestamp 1751429576
transform -1 0 36 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_81
timestamp 1751429576
transform -1 0 68 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_11
timestamp 1751429576
transform -1 0 92 0 1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_78
timestamp 1751429576
transform -1 0 124 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_10
timestamp 1751429576
transform -1 0 148 0 1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_82
timestamp 1751429576
transform 1 0 148 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_112
timestamp 1751429576
transform -1 0 212 0 1 1105
box -2 -3 34 103
use INVX2  INVX2_19
timestamp 1751429576
transform -1 0 228 0 1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_75
timestamp 1751429576
transform 1 0 228 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_102
timestamp 1751429576
transform 1 0 260 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_60
timestamp 1751429576
transform 1 0 292 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_57
timestamp 1751429576
transform -1 0 356 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_62
timestamp 1751429576
transform 1 0 356 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_104
timestamp 1751429576
transform -1 0 420 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_58
timestamp 1751429576
transform 1 0 420 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_53
timestamp 1751429576
transform -1 0 484 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_0_0
timestamp 1751429576
transform -1 0 492 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1751429576
transform -1 0 500 0 1 1105
box -2 -3 10 103
use INVX1  INVX1_33
timestamp 1751429576
transform -1 0 516 0 1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_49
timestamp 1751429576
transform 1 0 516 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_53
timestamp 1751429576
transform -1 0 564 0 1 1105
box -2 -3 26 103
use OR2X2  OR2X2_8
timestamp 1751429576
transform 1 0 564 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_42
timestamp 1751429576
transform -1 0 628 0 1 1105
box -2 -3 34 103
use INVX2  INVX2_14
timestamp 1751429576
transform -1 0 644 0 1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_34
timestamp 1751429576
transform -1 0 676 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_34
timestamp 1751429576
transform 1 0 676 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_70
timestamp 1751429576
transform 1 0 708 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_35
timestamp 1751429576
transform -1 0 772 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_28
timestamp 1751429576
transform 1 0 772 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_69
timestamp 1751429576
transform 1 0 788 0 1 1105
box -2 -3 34 103
use DFFSR  DFFSR_8
timestamp 1751429576
transform 1 0 820 0 1 1105
box -2 -3 178 103
use FILL  FILL_11_1_0
timestamp 1751429576
transform -1 0 1004 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1751429576
transform -1 0 1012 0 1 1105
box -2 -3 10 103
use NOR2X1  NOR2X1_18
timestamp 1751429576
transform -1 0 1036 0 1 1105
box -2 -3 26 103
use INVX2  INVX2_13
timestamp 1751429576
transform 1 0 1036 0 1 1105
box -2 -3 18 103
use AOI22X1  AOI22X1_7
timestamp 1751429576
transform -1 0 1092 0 1 1105
box -2 -3 42 103
use NAND3X1  NAND3X1_27
timestamp 1751429576
transform -1 0 1124 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_11
timestamp 1751429576
transform -1 0 1140 0 1 1105
box -2 -3 18 103
use AOI22X1  AOI22X1_9
timestamp 1751429576
transform 1 0 1140 0 1 1105
box -2 -3 42 103
use AOI22X1  AOI22X1_5
timestamp 1751429576
transform 1 0 1180 0 1 1105
box -2 -3 42 103
use DFFSR  DFFSR_4
timestamp 1751429576
transform 1 0 1220 0 1 1105
box -2 -3 178 103
use INVX1  INVX1_12
timestamp 1751429576
transform -1 0 1412 0 1 1105
box -2 -3 18 103
use BUFX2  BUFX2_5
timestamp 1751429576
transform 1 0 1412 0 1 1105
box -2 -3 26 103
use BUFX2  BUFX2_4
timestamp 1751429576
transform 1 0 1436 0 1 1105
box -2 -3 26 103
use BUFX2  BUFX2_9
timestamp 1751429576
transform 1 0 1460 0 1 1105
box -2 -3 26 103
use FILL  FILL_12_1
timestamp 1751429576
transform 1 0 1484 0 1 1105
box -2 -3 10 103
use FILL  FILL_12_2
timestamp 1751429576
transform 1 0 1492 0 1 1105
box -2 -3 10 103
use FILL  FILL_12_3
timestamp 1751429576
transform 1 0 1500 0 1 1105
box -2 -3 10 103
use NAND3X1  NAND3X1_84
timestamp 1751429576
transform -1 0 36 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_78
timestamp 1751429576
transform 1 0 36 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_18
timestamp 1751429576
transform -1 0 100 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_85
timestamp 1751429576
transform 1 0 100 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_126
timestamp 1751429576
transform 1 0 132 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_86
timestamp 1751429576
transform -1 0 196 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_11
timestamp 1751429576
transform 1 0 196 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_83
timestamp 1751429576
transform 1 0 228 0 -1 1305
box -2 -3 34 103
use AOI22X1  AOI22X1_11
timestamp 1751429576
transform -1 0 300 0 -1 1305
box -2 -3 42 103
use NOR2X1  NOR2X1_72
timestamp 1751429576
transform -1 0 324 0 -1 1305
box -2 -3 26 103
use NOR3X1  NOR3X1_6
timestamp 1751429576
transform 1 0 324 0 -1 1305
box -2 -3 66 103
use NAND3X1  NAND3X1_63
timestamp 1751429576
transform -1 0 420 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_103
timestamp 1751429576
transform 1 0 420 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_79
timestamp 1751429576
transform 1 0 452 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_0_0
timestamp 1751429576
transform 1 0 484 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1751429576
transform 1 0 492 0 -1 1305
box -2 -3 10 103
use NAND3X1  NAND3X1_61
timestamp 1751429576
transform 1 0 500 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_64
timestamp 1751429576
transform -1 0 564 0 -1 1305
box -2 -3 34 103
use NOR3X1  NOR3X1_5
timestamp 1751429576
transform -1 0 628 0 -1 1305
box -2 -3 66 103
use OAI21X1  OAI21X1_84
timestamp 1751429576
transform 1 0 628 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_34
timestamp 1751429576
transform 1 0 660 0 -1 1305
box -2 -3 18 103
use NAND3X1  NAND3X1_41
timestamp 1751429576
transform 1 0 676 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_32
timestamp 1751429576
transform -1 0 724 0 -1 1305
box -2 -3 18 103
use NAND3X1  NAND3X1_42
timestamp 1751429576
transform -1 0 756 0 -1 1305
box -2 -3 34 103
use INVX8  INVX8_1
timestamp 1751429576
transform -1 0 796 0 -1 1305
box -2 -3 42 103
use NAND3X1  NAND3X1_36
timestamp 1751429576
transform -1 0 828 0 -1 1305
box -2 -3 34 103
use DFFSR  DFFSR_7
timestamp 1751429576
transform 1 0 828 0 -1 1305
box -2 -3 178 103
use FILL  FILL_12_1_0
timestamp 1751429576
transform 1 0 1004 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1751429576
transform 1 0 1012 0 -1 1305
box -2 -3 10 103
use DFFSR  DFFSR_5
timestamp 1751429576
transform 1 0 1020 0 -1 1305
box -2 -3 178 103
use INVX1  INVX1_10
timestamp 1751429576
transform -1 0 1212 0 -1 1305
box -2 -3 18 103
use DFFSR  DFFSR_6
timestamp 1751429576
transform 1 0 1212 0 -1 1305
box -2 -3 178 103
use BUFX2  BUFX2_6
timestamp 1751429576
transform 1 0 1388 0 -1 1305
box -2 -3 26 103
use BUFX2  BUFX2_7
timestamp 1751429576
transform 1 0 1412 0 -1 1305
box -2 -3 26 103
use BUFX2  BUFX2_8
timestamp 1751429576
transform 1 0 1436 0 -1 1305
box -2 -3 26 103
use INVX2  INVX2_5
timestamp 1751429576
transform 1 0 1460 0 -1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_19
timestamp 1751429576
transform -1 0 1500 0 -1 1305
box -2 -3 26 103
use FILL  FILL_13_1
timestamp 1751429576
transform -1 0 1508 0 -1 1305
box -2 -3 10 103
<< labels >>
flabel metal6 s 480 -30 496 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 1000 -30 1016 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 574 -22 578 -18 7 FreeSans 24 270 0 0 a[0]
port 2 nsew
flabel metal3 s 1534 558 1538 562 3 FreeSans 24 0 0 0 a[1]
port 3 nsew
flabel metal3 s -26 668 -22 672 7 FreeSans 24 0 0 0 a[2]
port 4 nsew
flabel metal3 s -26 268 -22 272 7 FreeSans 24 0 0 0 a[3]
port 5 nsew
flabel metal2 s 782 -22 786 -18 7 FreeSans 24 270 0 0 a[4]
port 6 nsew
flabel metal2 s 518 -22 522 -18 7 FreeSans 24 270 0 0 a[5]
port 7 nsew
flabel metal2 s 702 -22 706 -18 7 FreeSans 24 270 0 0 a[6]
port 8 nsew
flabel metal2 s 662 -22 666 -18 7 FreeSans 24 270 0 0 a[7]
port 9 nsew
flabel metal2 s 638 -22 642 -18 7 FreeSans 24 270 0 0 b[0]
port 10 nsew
flabel metal2 s 430 -22 434 -18 7 FreeSans 24 270 0 0 b[1]
port 11 nsew
flabel metal2 s 542 -22 546 -18 7 FreeSans 24 270 0 0 b[2]
port 12 nsew
flabel metal2 s 270 -22 274 -18 7 FreeSans 24 270 0 0 b[3]
port 13 nsew
flabel metal2 s 806 -22 810 -18 7 FreeSans 24 270 0 0 b[4]
port 14 nsew
flabel metal2 s 678 -22 682 -18 7 FreeSans 24 270 0 0 b[5]
port 15 nsew
flabel metal2 s 750 -22 754 -18 7 FreeSans 24 270 0 0 b[6]
port 16 nsew
flabel metal2 s 1262 -22 1266 -18 7 FreeSans 24 270 0 0 b[7]
port 17 nsew
flabel metal2 s 910 1328 914 1332 3 FreeSans 24 90 0 0 clk
port 18 nsew
flabel metal2 s 774 1328 778 1332 3 FreeSans 24 90 0 0 rst
port 19 nsew
flabel metal2 s 1206 -22 1210 -18 7 FreeSans 24 270 0 0 en
port 20 nsew
flabel metal3 s 1534 1318 1538 1322 3 FreeSans 24 90 0 0 opcode[0]
port 21 nsew
flabel metal3 s 1534 278 1538 282 3 FreeSans 24 0 0 0 opcode[1]
port 22 nsew
flabel metal3 s 1534 258 1538 262 3 FreeSans 24 0 0 0 opcode[2]
port 23 nsew
flabel metal3 s 1534 848 1538 852 3 FreeSans 24 0 0 0 out[0]
port 24 nsew
flabel metal3 s 1534 948 1538 952 3 FreeSans 24 0 0 0 out[1]
port 25 nsew
flabel metal3 s 1534 968 1538 972 3 FreeSans 24 0 0 0 out[2]
port 26 nsew
flabel metal3 s 1534 1148 1538 1152 3 FreeSans 24 0 0 0 out[3]
port 27 nsew
flabel metal3 s 1534 1168 1538 1172 3 FreeSans 24 0 0 0 out[4]
port 28 nsew
flabel metal3 s 1534 1238 1538 1242 3 FreeSans 24 90 0 0 out[5]
port 29 nsew
flabel metal3 s 1534 1258 1538 1262 3 FreeSans 24 90 0 0 out[6]
port 30 nsew
flabel metal3 s 1534 1278 1538 1282 3 FreeSans 24 90 0 0 out[7]
port 31 nsew
flabel metal3 s 1534 1298 1538 1302 3 FreeSans 24 90 0 0 zero
port 32 nsew
<< end >>
